//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for physical tile: bram]
//	Author: Xifan TANG
//	Organization: University of Utah
//-------------------------------------------
//----- Time scale -----
`timescale 1ns / 1ps

// ----- BEGIN Grid Verilog module: grid_bram -----
//----- Default net type -----
`default_nettype wire

// ----- Verilog module for grid_bram -----
module grid_bram(scan_mode,
                 scan_enable,
                 global_reset,
                 rwm,
                 config_enable,
                 prog_clock,
                 top_width_0_height_0_subtile_0__pin_I00_0_,
                 top_width_0_height_0_subtile_0__pin_I00_1_,
                 top_width_0_height_0_subtile_0__pin_I00_2_,
                 top_width_0_height_0_subtile_0__pin_I00_3_,
                 top_width_0_height_0_subtile_0__pin_I00_4_,
                 top_width_0_height_0_subtile_0__pin_I00_5_,
                 top_width_0_height_0_subtile_0__pin_I00_6_,
                 top_width_0_height_0_subtile_0__pin_I00_7_,
                 top_width_0_height_0_subtile_0__pin_I00_8_,
                 top_width_0_height_0_subtile_0__pin_I00_9_,
                 top_width_0_height_0_subtile_0__pin_I00_10_,
                 top_width_0_height_0_subtile_0__pin_I00_11_,
                 top_width_0_height_0_subtile_0__pin_I10_0_,
                 top_width_0_height_0_subtile_0__pin_I10_1_,
                 top_width_0_height_0_subtile_0__pin_I10_2_,
                 top_width_0_height_0_subtile_0__pin_I10_3_,
                 top_width_0_height_0_subtile_0__pin_I10_4_,
                 top_width_0_height_0_subtile_0__pin_I10_5_,
                 top_width_0_height_0_subtile_0__pin_I10_6_,
                 top_width_0_height_0_subtile_0__pin_I10_7_,
                 top_width_0_height_0_subtile_0__pin_I10_8_,
                 top_width_0_height_0_subtile_0__pin_I10_9_,
                 top_width_0_height_0_subtile_0__pin_I10_10_,
                 top_width_0_height_0_subtile_0__pin_I10_11_,
                 top_width_0_height_0_subtile_0__pin_IS0_0_,
                 top_width_0_height_0_subtile_0__pin_IS0_1_,
                 top_width_0_height_0_subtile_0__pin_IS0_2_,
                 top_width_0_height_1_subtile_0__pin_I01_0_,
                 top_width_0_height_1_subtile_0__pin_I01_1_,
                 top_width_0_height_1_subtile_0__pin_I01_2_,
                 top_width_0_height_1_subtile_0__pin_I01_3_,
                 top_width_0_height_1_subtile_0__pin_I01_4_,
                 top_width_0_height_1_subtile_0__pin_I01_5_,
                 top_width_0_height_1_subtile_0__pin_I01_6_,
                 top_width_0_height_1_subtile_0__pin_I01_7_,
                 top_width_0_height_1_subtile_0__pin_I01_8_,
                 top_width_0_height_1_subtile_0__pin_I01_9_,
                 top_width_0_height_1_subtile_0__pin_I01_10_,
                 top_width_0_height_1_subtile_0__pin_I01_11_,
                 top_width_0_height_1_subtile_0__pin_I11_0_,
                 top_width_0_height_1_subtile_0__pin_I11_1_,
                 top_width_0_height_1_subtile_0__pin_I11_2_,
                 top_width_0_height_1_subtile_0__pin_I11_3_,
                 top_width_0_height_1_subtile_0__pin_I11_4_,
                 top_width_0_height_1_subtile_0__pin_I11_5_,
                 top_width_0_height_1_subtile_0__pin_I11_6_,
                 top_width_0_height_1_subtile_0__pin_I11_7_,
                 top_width_0_height_1_subtile_0__pin_I11_8_,
                 top_width_0_height_1_subtile_0__pin_I11_9_,
                 top_width_0_height_1_subtile_0__pin_I11_10_,
                 top_width_0_height_1_subtile_0__pin_I11_11_,
                 top_width_0_height_1_subtile_0__pin_IS1_0_,
                 top_width_0_height_1_subtile_0__pin_IS1_1_,
                 top_width_0_height_1_subtile_0__pin_IS1_2_,
                 top_width_0_height_2_subtile_0__pin_I02_0_,
                 top_width_0_height_2_subtile_0__pin_I02_1_,
                 top_width_0_height_2_subtile_0__pin_I02_2_,
                 top_width_0_height_2_subtile_0__pin_I02_3_,
                 top_width_0_height_2_subtile_0__pin_I02_4_,
                 top_width_0_height_2_subtile_0__pin_I02_5_,
                 top_width_0_height_2_subtile_0__pin_I02_6_,
                 top_width_0_height_2_subtile_0__pin_I02_7_,
                 top_width_0_height_2_subtile_0__pin_I02_8_,
                 top_width_0_height_2_subtile_0__pin_I02_9_,
                 top_width_0_height_2_subtile_0__pin_I02_10_,
                 top_width_0_height_2_subtile_0__pin_I02_11_,
                 top_width_0_height_2_subtile_0__pin_I12_0_,
                 top_width_0_height_2_subtile_0__pin_I12_1_,
                 top_width_0_height_2_subtile_0__pin_I12_2_,
                 top_width_0_height_2_subtile_0__pin_I12_3_,
                 top_width_0_height_2_subtile_0__pin_I12_4_,
                 top_width_0_height_2_subtile_0__pin_I12_5_,
                 top_width_0_height_2_subtile_0__pin_I12_6_,
                 top_width_0_height_2_subtile_0__pin_I12_7_,
                 top_width_0_height_2_subtile_0__pin_I12_8_,
                 top_width_0_height_2_subtile_0__pin_I12_9_,
                 top_width_0_height_2_subtile_0__pin_I12_10_,
                 top_width_0_height_2_subtile_0__pin_I12_11_,
                 top_width_0_height_2_subtile_0__pin_IS2_0_,
                 top_width_0_height_2_subtile_0__pin_IS2_1_,
                 top_width_0_height_2_subtile_0__pin_IS2_2_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_0_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_1_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_2_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_3_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_4_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_5_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_6_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_7_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_8_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_9_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_10_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_11_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_12_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_13_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_14_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_15_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_16_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_17_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_18_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_19_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_20_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_21_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_22_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_23_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_24_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_25_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_26_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_27_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_28_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_29_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_30_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_31_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_32_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_33_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_34_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_35_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_36_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_37_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_38_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_39_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_40_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_41_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_42_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_43_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_44_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_45_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_46_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_47_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_48_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_49_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_50_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_51_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_52_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_53_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_54_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_55_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_56_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_57_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_58_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_59_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_60_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_61_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_62_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_63_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_64_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_65_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_66_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_67_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_68_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_69_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_70_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_71_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_72_,
                 top_width_0_height_2_subtile_0__pin_PL_IN_73_,
                 right_width_0_height_0_subtile_0__pin_I20_0_,
                 right_width_0_height_0_subtile_0__pin_I20_1_,
                 right_width_0_height_0_subtile_0__pin_I20_2_,
                 right_width_0_height_0_subtile_0__pin_I20_3_,
                 right_width_0_height_0_subtile_0__pin_I20_4_,
                 right_width_0_height_0_subtile_0__pin_I20_5_,
                 right_width_0_height_0_subtile_0__pin_I20_6_,
                 right_width_0_height_0_subtile_0__pin_I20_7_,
                 right_width_0_height_0_subtile_0__pin_I20_8_,
                 right_width_0_height_0_subtile_0__pin_I20_9_,
                 right_width_0_height_0_subtile_0__pin_I20_10_,
                 right_width_0_height_0_subtile_0__pin_I20_11_,
                 right_width_0_height_0_subtile_0__pin_I30_0_,
                 right_width_0_height_0_subtile_0__pin_I30_1_,
                 right_width_0_height_0_subtile_0__pin_I30_2_,
                 right_width_0_height_0_subtile_0__pin_I30_3_,
                 right_width_0_height_0_subtile_0__pin_I30_4_,
                 right_width_0_height_0_subtile_0__pin_I30_5_,
                 right_width_0_height_0_subtile_0__pin_I30_6_,
                 right_width_0_height_0_subtile_0__pin_I30_7_,
                 right_width_0_height_0_subtile_0__pin_I30_8_,
                 right_width_0_height_0_subtile_0__pin_I30_9_,
                 right_width_0_height_0_subtile_0__pin_I30_10_,
                 right_width_0_height_0_subtile_0__pin_I30_11_,
                 right_width_0_height_0_subtile_0__pin_IS0_3_,
                 right_width_0_height_0_subtile_0__pin_IS0_4_,
                 right_width_0_height_0_subtile_0__pin_IS0_5_,
                 right_width_0_height_1_subtile_0__pin_I21_0_,
                 right_width_0_height_1_subtile_0__pin_I21_1_,
                 right_width_0_height_1_subtile_0__pin_I21_2_,
                 right_width_0_height_1_subtile_0__pin_I21_3_,
                 right_width_0_height_1_subtile_0__pin_I21_4_,
                 right_width_0_height_1_subtile_0__pin_I21_5_,
                 right_width_0_height_1_subtile_0__pin_I21_6_,
                 right_width_0_height_1_subtile_0__pin_I21_7_,
                 right_width_0_height_1_subtile_0__pin_I21_8_,
                 right_width_0_height_1_subtile_0__pin_I21_9_,
                 right_width_0_height_1_subtile_0__pin_I21_10_,
                 right_width_0_height_1_subtile_0__pin_I21_11_,
                 right_width_0_height_1_subtile_0__pin_I31_0_,
                 right_width_0_height_1_subtile_0__pin_I31_1_,
                 right_width_0_height_1_subtile_0__pin_I31_2_,
                 right_width_0_height_1_subtile_0__pin_I31_3_,
                 right_width_0_height_1_subtile_0__pin_I31_4_,
                 right_width_0_height_1_subtile_0__pin_I31_5_,
                 right_width_0_height_1_subtile_0__pin_I31_6_,
                 right_width_0_height_1_subtile_0__pin_I31_7_,
                 right_width_0_height_1_subtile_0__pin_I31_8_,
                 right_width_0_height_1_subtile_0__pin_I31_9_,
                 right_width_0_height_1_subtile_0__pin_I31_10_,
                 right_width_0_height_1_subtile_0__pin_I31_11_,
                 right_width_0_height_1_subtile_0__pin_IS1_3_,
                 right_width_0_height_1_subtile_0__pin_IS1_4_,
                 right_width_0_height_1_subtile_0__pin_IS1_5_,
                 right_width_0_height_2_subtile_0__pin_I22_0_,
                 right_width_0_height_2_subtile_0__pin_I22_1_,
                 right_width_0_height_2_subtile_0__pin_I22_2_,
                 right_width_0_height_2_subtile_0__pin_I22_3_,
                 right_width_0_height_2_subtile_0__pin_I22_4_,
                 right_width_0_height_2_subtile_0__pin_I22_5_,
                 right_width_0_height_2_subtile_0__pin_I22_6_,
                 right_width_0_height_2_subtile_0__pin_I22_7_,
                 right_width_0_height_2_subtile_0__pin_I22_8_,
                 right_width_0_height_2_subtile_0__pin_I22_9_,
                 right_width_0_height_2_subtile_0__pin_I22_10_,
                 right_width_0_height_2_subtile_0__pin_I22_11_,
                 right_width_0_height_2_subtile_0__pin_I32_0_,
                 right_width_0_height_2_subtile_0__pin_I32_1_,
                 right_width_0_height_2_subtile_0__pin_I32_2_,
                 right_width_0_height_2_subtile_0__pin_I32_3_,
                 right_width_0_height_2_subtile_0__pin_I32_4_,
                 right_width_0_height_2_subtile_0__pin_I32_5_,
                 right_width_0_height_2_subtile_0__pin_I32_6_,
                 right_width_0_height_2_subtile_0__pin_I32_7_,
                 right_width_0_height_2_subtile_0__pin_I32_8_,
                 right_width_0_height_2_subtile_0__pin_I32_9_,
                 right_width_0_height_2_subtile_0__pin_I32_10_,
                 right_width_0_height_2_subtile_0__pin_I32_11_,
                 right_width_0_height_2_subtile_0__pin_IS2_3_,
                 right_width_0_height_2_subtile_0__pin_IS2_4_,
                 right_width_0_height_2_subtile_0__pin_IS2_5_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_0_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_1_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_2_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_3_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_4_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_5_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_6_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_7_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_8_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_9_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_10_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_11_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_12_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_13_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_14_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_15_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_16_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_17_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_18_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_19_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_20_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_21_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_22_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_23_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_24_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_25_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_26_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_27_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_28_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_29_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_30_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_31_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_32_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_33_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_34_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_35_,
                 left_width_0_height_0_subtile_0__pin_sc_in_0_,
                 left_width_0_height_0_subtile_0__pin_sc_in_1_,
                 left_width_0_height_0_subtile_0__pin_sc_in_2_,
                 left_width_0_height_0_subtile_0__pin_sc_in_3_,
                 left_width_0_height_0_subtile_0__pin_sc_in_4_,
                 left_width_0_height_0_subtile_0__pin_sc_in_5_,
                 left_width_0_height_0_subtile_0__pin_sc_in_6_,
                 left_width_0_height_0_subtile_0__pin_sc_in_7_,
                 left_width_0_height_0_subtile_0__pin_sc_in_8_,
                 left_width_0_height_0_subtile_0__pin_sc_in_9_,
                 left_width_0_height_0_subtile_0__pin_sc_in_10_,
                 left_width_0_height_0_subtile_0__pin_sc_in_11_,
                 left_width_0_height_0_subtile_0__pin_sc_in_12_,
                 left_width_0_height_0_subtile_0__pin_sc_in_13_,
                 left_width_0_height_0_subtile_0__pin_sc_in_14_,
                 left_width_0_height_0_subtile_0__pin_sc_in_15_,
                 left_width_0_height_0_subtile_0__pin_sc_in_16_,
                 left_width_0_height_0_subtile_0__pin_sc_in_17_,
                 left_width_0_height_0_subtile_0__pin_sc_in_18_,
                 left_width_0_height_0_subtile_0__pin_sc_in_19_,
                 left_width_0_height_0_subtile_0__pin_sc_in_20_,
                 left_width_0_height_0_subtile_0__pin_sc_in_21_,
                 left_width_0_height_0_subtile_0__pin_sc_in_22_,
                 left_width_0_height_0_subtile_0__pin_sc_in_23_,
                 left_width_0_height_0_subtile_0__pin_sc_in_24_,
                 left_width_0_height_0_subtile_0__pin_sc_in_25_,
                 left_width_0_height_0_subtile_0__pin_sc_in_26_,
                 left_width_0_height_0_subtile_0__pin_sc_in_27_,
                 left_width_0_height_0_subtile_0__pin_sc_in_28_,
                 left_width_0_height_0_subtile_0__pin_sc_in_29_,
                 left_width_0_height_0_subtile_0__pin_sc_in_30_,
                 left_width_0_height_0_subtile_0__pin_sc_in_31_,
                 left_width_0_height_0_subtile_0__pin_sc_in_32_,
                 left_width_0_height_0_subtile_0__pin_sc_in_33_,
                 left_width_0_height_0_subtile_0__pin_sc_in_34_,
                 left_width_0_height_0_subtile_0__pin_sc_in_35_,
                 left_width_0_height_0_subtile_0__pin_sc_in_36_,
                 left_width_0_height_0_subtile_0__pin_sc_in_37_,
                 left_width_0_height_0_subtile_0__pin_sc_in_38_,
                 left_width_0_height_0_subtile_0__pin_sc_in_39_,
                 left_width_0_height_0_subtile_0__pin_sc_in_40_,
                 left_width_0_height_0_subtile_0__pin_sc_in_41_,
                 left_width_0_height_0_subtile_0__pin_sc_in_42_,
                 left_width_0_height_0_subtile_0__pin_sc_in_43_,
                 left_width_0_height_0_subtile_0__pin_sc_in_44_,
                 left_width_0_height_0_subtile_0__pin_sc_in_45_,
                 left_width_0_height_0_subtile_0__pin_sc_in_46_,
                 left_width_0_height_0_subtile_0__pin_sc_in_47_,
                 left_width_0_height_0_subtile_0__pin_clk_0_,
                 left_width_0_height_0_subtile_0__pin_clk_1_,
                 left_width_0_height_0_subtile_0__pin_clk_2_,
                 left_width_0_height_0_subtile_0__pin_clk_3_,
                 left_width_0_height_0_subtile_0__pin_clk_4_,
                 left_width_0_height_0_subtile_0__pin_clk_5_,
                 left_width_0_height_0_subtile_0__pin_clk_6_,
                 left_width_0_height_0_subtile_0__pin_clk_7_,
                 left_width_0_height_0_subtile_0__pin_clk_8_,
                 left_width_0_height_0_subtile_0__pin_clk_9_,
                 left_width_0_height_0_subtile_0__pin_clk_10_,
                 left_width_0_height_0_subtile_0__pin_clk_11_,
                 left_width_0_height_0_subtile_0__pin_clk_12_,
                 left_width_0_height_0_subtile_0__pin_clk_13_,
                 left_width_0_height_0_subtile_0__pin_clk_14_,
                 left_width_0_height_0_subtile_0__pin_clk_15_,
                 left_width_0_height_1_subtile_0__pin_RAM_ID_i_0_,
                 left_width_0_height_1_subtile_0__pin_RAM_ID_i_1_,
                 left_width_0_height_1_subtile_0__pin_RAM_ID_i_2_,
                 left_width_0_height_1_subtile_0__pin_RAM_ID_i_3_,
                 left_width_0_height_1_subtile_0__pin_RAM_ID_i_4_,
                 left_width_0_height_1_subtile_0__pin_RAM_ID_i_5_,
                 left_width_0_height_1_subtile_0__pin_RAM_ID_i_6_,
                 left_width_0_height_1_subtile_0__pin_RAM_ID_i_7_,
                 left_width_0_height_1_subtile_0__pin_RAM_ID_i_8_,
                 left_width_0_height_1_subtile_0__pin_RAM_ID_i_9_,
                 left_width_0_height_1_subtile_0__pin_RAM_ID_i_10_,
                 left_width_0_height_1_subtile_0__pin_RAM_ID_i_11_,
                 left_width_0_height_1_subtile_0__pin_RAM_ID_i_12_,
                 left_width_0_height_1_subtile_0__pin_RAM_ID_i_13_,
                 left_width_0_height_1_subtile_0__pin_RAM_ID_i_14_,
                 left_width_0_height_1_subtile_0__pin_RAM_ID_i_15_,
                 left_width_0_height_1_subtile_0__pin_RAM_ID_i_16_,
                 left_width_0_height_1_subtile_0__pin_RAM_ID_i_17_,
                 left_width_0_height_1_subtile_0__pin_RAM_ID_i_18_,
                 left_width_0_height_1_subtile_0__pin_RAM_ID_i_19_,
                 ccff_head,
                 top_width_0_height_0_subtile_0__pin_O0_0_,
                 top_width_0_height_0_subtile_0__pin_O0_1_,
                 top_width_0_height_0_subtile_0__pin_O0_2_,
                 top_width_0_height_0_subtile_0__pin_O0_3_,
                 top_width_0_height_0_subtile_0__pin_O0_4_,
                 top_width_0_height_0_subtile_0__pin_O0_5_,
                 top_width_0_height_0_subtile_0__pin_O0_6_,
                 top_width_0_height_0_subtile_0__pin_O0_7_,
                 top_width_0_height_0_subtile_0__pin_O0_8_,
                 top_width_0_height_0_subtile_0__pin_O0_9_,
                 top_width_0_height_0_subtile_0__pin_O0_10_,
                 top_width_0_height_0_subtile_0__pin_O0_11_,
                 top_width_0_height_1_subtile_0__pin_O1_0_,
                 top_width_0_height_1_subtile_0__pin_O1_1_,
                 top_width_0_height_1_subtile_0__pin_O1_2_,
                 top_width_0_height_1_subtile_0__pin_O1_3_,
                 top_width_0_height_1_subtile_0__pin_O1_4_,
                 top_width_0_height_1_subtile_0__pin_O1_5_,
                 top_width_0_height_1_subtile_0__pin_O1_6_,
                 top_width_0_height_1_subtile_0__pin_O1_7_,
                 top_width_0_height_1_subtile_0__pin_O1_8_,
                 top_width_0_height_1_subtile_0__pin_O1_9_,
                 top_width_0_height_1_subtile_0__pin_O1_10_,
                 top_width_0_height_1_subtile_0__pin_O1_11_,
                 top_width_0_height_2_subtile_0__pin_O2_0_,
                 top_width_0_height_2_subtile_0__pin_O2_1_,
                 top_width_0_height_2_subtile_0__pin_O2_2_,
                 top_width_0_height_2_subtile_0__pin_O2_3_,
                 top_width_0_height_2_subtile_0__pin_O2_4_,
                 top_width_0_height_2_subtile_0__pin_O2_5_,
                 top_width_0_height_2_subtile_0__pin_O2_6_,
                 top_width_0_height_2_subtile_0__pin_O2_7_,
                 top_width_0_height_2_subtile_0__pin_O2_8_,
                 top_width_0_height_2_subtile_0__pin_O2_9_,
                 top_width_0_height_2_subtile_0__pin_O2_10_,
                 top_width_0_height_2_subtile_0__pin_O2_11_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_0_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_1_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_2_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_3_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_4_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_5_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_6_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_7_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_8_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_9_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_10_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_11_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_12_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_13_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_14_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_15_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_16_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_17_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_18_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_19_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_20_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_21_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_22_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_23_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_24_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_25_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_26_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_27_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_28_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_29_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_30_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_31_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_32_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_33_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_34_,
                 top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_35_,
                 right_width_0_height_0_subtile_0__pin_O0_12_,
                 right_width_0_height_0_subtile_0__pin_O0_13_,
                 right_width_0_height_0_subtile_0__pin_O0_14_,
                 right_width_0_height_0_subtile_0__pin_O0_15_,
                 right_width_0_height_0_subtile_0__pin_O0_16_,
                 right_width_0_height_0_subtile_0__pin_O0_17_,
                 right_width_0_height_0_subtile_0__pin_O0_18_,
                 right_width_0_height_0_subtile_0__pin_O0_19_,
                 right_width_0_height_0_subtile_0__pin_O0_20_,
                 right_width_0_height_0_subtile_0__pin_O0_21_,
                 right_width_0_height_0_subtile_0__pin_O0_22_,
                 right_width_0_height_0_subtile_0__pin_O0_23_,
                 right_width_0_height_0_subtile_0__pin_sc_out_0_,
                 right_width_0_height_0_subtile_0__pin_sc_out_1_,
                 right_width_0_height_0_subtile_0__pin_sc_out_2_,
                 right_width_0_height_0_subtile_0__pin_sc_out_3_,
                 right_width_0_height_0_subtile_0__pin_sc_out_4_,
                 right_width_0_height_0_subtile_0__pin_sc_out_5_,
                 right_width_0_height_0_subtile_0__pin_sc_out_6_,
                 right_width_0_height_0_subtile_0__pin_sc_out_7_,
                 right_width_0_height_0_subtile_0__pin_sc_out_8_,
                 right_width_0_height_0_subtile_0__pin_sc_out_9_,
                 right_width_0_height_0_subtile_0__pin_sc_out_10_,
                 right_width_0_height_0_subtile_0__pin_sc_out_11_,
                 right_width_0_height_0_subtile_0__pin_sc_out_12_,
                 right_width_0_height_0_subtile_0__pin_sc_out_13_,
                 right_width_0_height_0_subtile_0__pin_sc_out_14_,
                 right_width_0_height_0_subtile_0__pin_sc_out_15_,
                 right_width_0_height_0_subtile_0__pin_sc_out_16_,
                 right_width_0_height_0_subtile_0__pin_sc_out_17_,
                 right_width_0_height_0_subtile_0__pin_sc_out_18_,
                 right_width_0_height_0_subtile_0__pin_sc_out_19_,
                 right_width_0_height_0_subtile_0__pin_sc_out_20_,
                 right_width_0_height_0_subtile_0__pin_sc_out_21_,
                 right_width_0_height_0_subtile_0__pin_sc_out_22_,
                 right_width_0_height_0_subtile_0__pin_sc_out_23_,
                 right_width_0_height_0_subtile_0__pin_sc_out_24_,
                 right_width_0_height_0_subtile_0__pin_sc_out_25_,
                 right_width_0_height_0_subtile_0__pin_sc_out_26_,
                 right_width_0_height_0_subtile_0__pin_sc_out_27_,
                 right_width_0_height_0_subtile_0__pin_sc_out_28_,
                 right_width_0_height_0_subtile_0__pin_sc_out_29_,
                 right_width_0_height_0_subtile_0__pin_sc_out_30_,
                 right_width_0_height_0_subtile_0__pin_sc_out_31_,
                 right_width_0_height_0_subtile_0__pin_sc_out_32_,
                 right_width_0_height_0_subtile_0__pin_sc_out_33_,
                 right_width_0_height_0_subtile_0__pin_sc_out_34_,
                 right_width_0_height_0_subtile_0__pin_sc_out_35_,
                 right_width_0_height_0_subtile_0__pin_sc_out_36_,
                 right_width_0_height_0_subtile_0__pin_sc_out_37_,
                 right_width_0_height_0_subtile_0__pin_sc_out_38_,
                 right_width_0_height_0_subtile_0__pin_sc_out_39_,
                 right_width_0_height_0_subtile_0__pin_sc_out_40_,
                 right_width_0_height_0_subtile_0__pin_sc_out_41_,
                 right_width_0_height_0_subtile_0__pin_sc_out_42_,
                 right_width_0_height_0_subtile_0__pin_sc_out_43_,
                 right_width_0_height_0_subtile_0__pin_sc_out_44_,
                 right_width_0_height_0_subtile_0__pin_sc_out_45_,
                 right_width_0_height_0_subtile_0__pin_sc_out_46_,
                 right_width_0_height_0_subtile_0__pin_sc_out_47_,
                 right_width_0_height_1_subtile_0__pin_O1_12_,
                 right_width_0_height_1_subtile_0__pin_O1_13_,
                 right_width_0_height_1_subtile_0__pin_O1_14_,
                 right_width_0_height_1_subtile_0__pin_O1_15_,
                 right_width_0_height_1_subtile_0__pin_O1_16_,
                 right_width_0_height_1_subtile_0__pin_O1_17_,
                 right_width_0_height_1_subtile_0__pin_O1_18_,
                 right_width_0_height_1_subtile_0__pin_O1_19_,
                 right_width_0_height_1_subtile_0__pin_O1_20_,
                 right_width_0_height_1_subtile_0__pin_O1_21_,
                 right_width_0_height_1_subtile_0__pin_O1_22_,
                 right_width_0_height_1_subtile_0__pin_O1_23_,
                 right_width_0_height_2_subtile_0__pin_O2_12_,
                 right_width_0_height_2_subtile_0__pin_O2_13_,
                 right_width_0_height_2_subtile_0__pin_O2_14_,
                 right_width_0_height_2_subtile_0__pin_O2_15_,
                 right_width_0_height_2_subtile_0__pin_O2_16_,
                 right_width_0_height_2_subtile_0__pin_O2_17_,
                 right_width_0_height_2_subtile_0__pin_O2_18_,
                 right_width_0_height_2_subtile_0__pin_O2_19_,
                 right_width_0_height_2_subtile_0__pin_O2_20_,
                 right_width_0_height_2_subtile_0__pin_O2_21_,
                 right_width_0_height_2_subtile_0__pin_O2_22_,
                 right_width_0_height_2_subtile_0__pin_O2_23_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_0_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_1_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_2_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_3_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_4_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_5_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_6_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_7_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_8_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_9_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_10_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_11_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_12_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_13_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_14_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_15_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_16_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_17_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_18_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_19_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_20_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_21_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_22_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_23_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_24_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_25_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_26_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_27_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_28_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_29_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_30_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_31_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_32_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_33_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_34_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_35_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_36_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_37_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_38_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_39_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_40_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_41_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_42_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_43_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_44_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_45_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_46_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_47_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_48_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_49_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_50_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_51_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_52_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_53_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_54_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_55_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_56_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_57_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_58_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_59_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_60_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_61_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_62_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_63_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_64_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_65_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_66_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_67_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_68_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_69_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_70_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_71_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_72_,
                 bottom_width_0_height_0_subtile_0__pin_PL_OUT_73_,
                 ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] scan_mode;
//----- GLOBAL PORTS -----
input [0:0] scan_enable;
//----- GLOBAL PORTS -----
input [0:0] global_reset;
//----- GLOBAL PORTS -----
input [0:2] rwm;
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_clock;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I00_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I00_1_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I00_2_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I00_3_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I00_4_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I00_5_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I00_6_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I00_7_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I00_8_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I00_9_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I00_10_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I00_11_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I10_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I10_1_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I10_2_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I10_3_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I10_4_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I10_5_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I10_6_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I10_7_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I10_8_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I10_9_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I10_10_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I10_11_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_IS0_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_IS0_1_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_IS0_2_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I01_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I01_1_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I01_2_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I01_3_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I01_4_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I01_5_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I01_6_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I01_7_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I01_8_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I01_9_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I01_10_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I01_11_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I11_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I11_1_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I11_2_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I11_3_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I11_4_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I11_5_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I11_6_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I11_7_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I11_8_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I11_9_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I11_10_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I11_11_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_IS1_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_IS1_1_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_IS1_2_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I02_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I02_1_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I02_2_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I02_3_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I02_4_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I02_5_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I02_6_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I02_7_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I02_8_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I02_9_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I02_10_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I02_11_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I12_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I12_1_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I12_2_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I12_3_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I12_4_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I12_5_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I12_6_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I12_7_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I12_8_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I12_9_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I12_10_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I12_11_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_IS2_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_IS2_1_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_IS2_2_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_1_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_2_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_3_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_4_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_5_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_6_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_7_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_8_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_9_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_10_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_11_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_12_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_13_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_14_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_15_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_16_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_17_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_18_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_19_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_20_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_21_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_22_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_23_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_24_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_25_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_26_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_27_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_28_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_29_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_30_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_31_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_32_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_33_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_34_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_35_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_36_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_37_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_38_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_39_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_40_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_41_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_42_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_43_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_44_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_45_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_46_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_47_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_48_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_49_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_50_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_51_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_52_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_53_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_54_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_55_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_56_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_57_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_58_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_59_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_60_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_61_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_62_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_63_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_64_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_65_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_66_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_67_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_68_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_69_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_70_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_71_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_72_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_PL_IN_73_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I20_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I20_1_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I20_2_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I20_3_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I20_4_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I20_5_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I20_6_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I20_7_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I20_8_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I20_9_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I20_10_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I20_11_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I30_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I30_1_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I30_2_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I30_3_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I30_4_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I30_5_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I30_6_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I30_7_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I30_8_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I30_9_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I30_10_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I30_11_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_IS0_3_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_IS0_4_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_IS0_5_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I21_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I21_1_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I21_2_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I21_3_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I21_4_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I21_5_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I21_6_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I21_7_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I21_8_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I21_9_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I21_10_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I21_11_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I31_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I31_1_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I31_2_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I31_3_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I31_4_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I31_5_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I31_6_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I31_7_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I31_8_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I31_9_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I31_10_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I31_11_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_IS1_3_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_IS1_4_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_IS1_5_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I22_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I22_1_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I22_2_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I22_3_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I22_4_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I22_5_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I22_6_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I22_7_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I22_8_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I22_9_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I22_10_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I22_11_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I32_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I32_1_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I32_2_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I32_3_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I32_4_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I32_5_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I32_6_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I32_7_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I32_8_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I32_9_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I32_10_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I32_11_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_IS2_3_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_IS2_4_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_IS2_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_16_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_17_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_18_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_19_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_20_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_21_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_22_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_23_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_24_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_25_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_26_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_27_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_28_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_29_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_30_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_31_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_32_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_33_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_34_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_35_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_1_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_2_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_3_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_4_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_5_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_6_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_7_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_8_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_9_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_10_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_11_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_12_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_13_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_14_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_15_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_16_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_17_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_18_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_19_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_20_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_21_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_22_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_23_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_24_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_25_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_26_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_27_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_28_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_29_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_30_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_31_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_32_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_33_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_34_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_35_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_36_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_37_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_38_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_39_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_40_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_41_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_42_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_43_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_44_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_45_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_46_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_47_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_RAM_ID_i_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_RAM_ID_i_1_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_RAM_ID_i_2_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_RAM_ID_i_3_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_RAM_ID_i_4_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_RAM_ID_i_5_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_RAM_ID_i_6_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_RAM_ID_i_7_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_RAM_ID_i_8_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_RAM_ID_i_9_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_RAM_ID_i_10_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_RAM_ID_i_11_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_RAM_ID_i_12_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_RAM_ID_i_13_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_RAM_ID_i_14_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_RAM_ID_i_15_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_RAM_ID_i_16_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_RAM_ID_i_17_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_RAM_ID_i_18_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_1_subtile_0__pin_RAM_ID_i_19_;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_O0_0_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_O0_1_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_O0_2_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_O0_3_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_O0_4_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_O0_5_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_O0_6_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_O0_7_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_O0_8_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_O0_9_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_O0_10_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_O0_11_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_1_subtile_0__pin_O1_0_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_1_subtile_0__pin_O1_1_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_1_subtile_0__pin_O1_2_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_1_subtile_0__pin_O1_3_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_1_subtile_0__pin_O1_4_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_1_subtile_0__pin_O1_5_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_1_subtile_0__pin_O1_6_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_1_subtile_0__pin_O1_7_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_1_subtile_0__pin_O1_8_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_1_subtile_0__pin_O1_9_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_1_subtile_0__pin_O1_10_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_1_subtile_0__pin_O1_11_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_O2_0_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_O2_1_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_O2_2_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_O2_3_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_O2_4_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_O2_5_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_O2_6_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_O2_7_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_O2_8_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_O2_9_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_O2_10_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_O2_11_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_0_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_1_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_2_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_3_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_4_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_5_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_6_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_7_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_8_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_9_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_10_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_11_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_12_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_13_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_14_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_15_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_16_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_17_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_18_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_19_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_20_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_21_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_22_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_23_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_24_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_25_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_26_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_27_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_28_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_29_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_30_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_31_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_32_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_33_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_34_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_35_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_O0_12_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_O0_13_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_O0_14_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_O0_15_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_O0_16_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_O0_17_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_O0_18_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_O0_19_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_O0_20_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_O0_21_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_O0_22_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_O0_23_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_1_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_2_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_3_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_4_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_5_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_6_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_7_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_8_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_9_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_10_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_11_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_12_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_13_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_14_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_15_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_16_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_17_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_18_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_19_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_20_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_21_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_22_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_23_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_24_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_25_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_26_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_27_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_28_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_29_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_30_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_31_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_32_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_33_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_34_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_35_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_36_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_37_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_38_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_39_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_40_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_41_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_42_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_43_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_44_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_45_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_46_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_47_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_O1_12_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_O1_13_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_O1_14_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_O1_15_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_O1_16_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_O1_17_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_O1_18_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_O1_19_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_O1_20_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_O1_21_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_O1_22_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_O1_23_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_2_subtile_0__pin_O2_12_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_2_subtile_0__pin_O2_13_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_2_subtile_0__pin_O2_14_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_2_subtile_0__pin_O2_15_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_2_subtile_0__pin_O2_16_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_2_subtile_0__pin_O2_17_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_2_subtile_0__pin_O2_18_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_2_subtile_0__pin_O2_19_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_2_subtile_0__pin_O2_20_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_2_subtile_0__pin_O2_21_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_2_subtile_0__pin_O2_22_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_2_subtile_0__pin_O2_23_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_1_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_2_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_3_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_4_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_5_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_6_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_7_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_8_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_9_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_10_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_11_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_12_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_13_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_14_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_15_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_16_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_17_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_18_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_19_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_20_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_21_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_22_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_23_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_24_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_25_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_26_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_27_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_28_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_29_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_30_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_31_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_32_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_33_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_34_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_35_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_36_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_37_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_38_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_39_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_40_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_41_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_42_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_43_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_44_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_45_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_46_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_47_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_48_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_49_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_50_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_51_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_52_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_53_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_54_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_55_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_56_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_57_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_58_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_59_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_60_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_61_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_62_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_63_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_64_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_65_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_66_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_67_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_68_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_69_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_70_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_71_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_72_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_OUT_73_;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	logical_tile_bram_mode_bram_ logical_tile_bram_mode_bram__0 (
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.global_reset(global_reset),
		.rwm(rwm[0:2]),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.bram_I00({top_width_0_height_0_subtile_0__pin_I00_0_, top_width_0_height_0_subtile_0__pin_I00_1_, top_width_0_height_0_subtile_0__pin_I00_2_, top_width_0_height_0_subtile_0__pin_I00_3_, top_width_0_height_0_subtile_0__pin_I00_4_, top_width_0_height_0_subtile_0__pin_I00_5_, top_width_0_height_0_subtile_0__pin_I00_6_, top_width_0_height_0_subtile_0__pin_I00_7_, top_width_0_height_0_subtile_0__pin_I00_8_, top_width_0_height_0_subtile_0__pin_I00_9_, top_width_0_height_0_subtile_0__pin_I00_10_, top_width_0_height_0_subtile_0__pin_I00_11_}),
		.bram_I10({top_width_0_height_0_subtile_0__pin_I10_0_, top_width_0_height_0_subtile_0__pin_I10_1_, top_width_0_height_0_subtile_0__pin_I10_2_, top_width_0_height_0_subtile_0__pin_I10_3_, top_width_0_height_0_subtile_0__pin_I10_4_, top_width_0_height_0_subtile_0__pin_I10_5_, top_width_0_height_0_subtile_0__pin_I10_6_, top_width_0_height_0_subtile_0__pin_I10_7_, top_width_0_height_0_subtile_0__pin_I10_8_, top_width_0_height_0_subtile_0__pin_I10_9_, top_width_0_height_0_subtile_0__pin_I10_10_, top_width_0_height_0_subtile_0__pin_I10_11_}),
		.bram_I20({right_width_0_height_0_subtile_0__pin_I20_0_, right_width_0_height_0_subtile_0__pin_I20_1_, right_width_0_height_0_subtile_0__pin_I20_2_, right_width_0_height_0_subtile_0__pin_I20_3_, right_width_0_height_0_subtile_0__pin_I20_4_, right_width_0_height_0_subtile_0__pin_I20_5_, right_width_0_height_0_subtile_0__pin_I20_6_, right_width_0_height_0_subtile_0__pin_I20_7_, right_width_0_height_0_subtile_0__pin_I20_8_, right_width_0_height_0_subtile_0__pin_I20_9_, right_width_0_height_0_subtile_0__pin_I20_10_, right_width_0_height_0_subtile_0__pin_I20_11_}),
		.bram_I30({right_width_0_height_0_subtile_0__pin_I30_0_, right_width_0_height_0_subtile_0__pin_I30_1_, right_width_0_height_0_subtile_0__pin_I30_2_, right_width_0_height_0_subtile_0__pin_I30_3_, right_width_0_height_0_subtile_0__pin_I30_4_, right_width_0_height_0_subtile_0__pin_I30_5_, right_width_0_height_0_subtile_0__pin_I30_6_, right_width_0_height_0_subtile_0__pin_I30_7_, right_width_0_height_0_subtile_0__pin_I30_8_, right_width_0_height_0_subtile_0__pin_I30_9_, right_width_0_height_0_subtile_0__pin_I30_10_, right_width_0_height_0_subtile_0__pin_I30_11_}),
		.bram_IS0({top_width_0_height_0_subtile_0__pin_IS0_0_, top_width_0_height_0_subtile_0__pin_IS0_1_, top_width_0_height_0_subtile_0__pin_IS0_2_, right_width_0_height_0_subtile_0__pin_IS0_3_, right_width_0_height_0_subtile_0__pin_IS0_4_, right_width_0_height_0_subtile_0__pin_IS0_5_}),
		.bram_I01({top_width_0_height_1_subtile_0__pin_I01_0_, top_width_0_height_1_subtile_0__pin_I01_1_, top_width_0_height_1_subtile_0__pin_I01_2_, top_width_0_height_1_subtile_0__pin_I01_3_, top_width_0_height_1_subtile_0__pin_I01_4_, top_width_0_height_1_subtile_0__pin_I01_5_, top_width_0_height_1_subtile_0__pin_I01_6_, top_width_0_height_1_subtile_0__pin_I01_7_, top_width_0_height_1_subtile_0__pin_I01_8_, top_width_0_height_1_subtile_0__pin_I01_9_, top_width_0_height_1_subtile_0__pin_I01_10_, top_width_0_height_1_subtile_0__pin_I01_11_}),
		.bram_I11({top_width_0_height_1_subtile_0__pin_I11_0_, top_width_0_height_1_subtile_0__pin_I11_1_, top_width_0_height_1_subtile_0__pin_I11_2_, top_width_0_height_1_subtile_0__pin_I11_3_, top_width_0_height_1_subtile_0__pin_I11_4_, top_width_0_height_1_subtile_0__pin_I11_5_, top_width_0_height_1_subtile_0__pin_I11_6_, top_width_0_height_1_subtile_0__pin_I11_7_, top_width_0_height_1_subtile_0__pin_I11_8_, top_width_0_height_1_subtile_0__pin_I11_9_, top_width_0_height_1_subtile_0__pin_I11_10_, top_width_0_height_1_subtile_0__pin_I11_11_}),
		.bram_I21({right_width_0_height_1_subtile_0__pin_I21_0_, right_width_0_height_1_subtile_0__pin_I21_1_, right_width_0_height_1_subtile_0__pin_I21_2_, right_width_0_height_1_subtile_0__pin_I21_3_, right_width_0_height_1_subtile_0__pin_I21_4_, right_width_0_height_1_subtile_0__pin_I21_5_, right_width_0_height_1_subtile_0__pin_I21_6_, right_width_0_height_1_subtile_0__pin_I21_7_, right_width_0_height_1_subtile_0__pin_I21_8_, right_width_0_height_1_subtile_0__pin_I21_9_, right_width_0_height_1_subtile_0__pin_I21_10_, right_width_0_height_1_subtile_0__pin_I21_11_}),
		.bram_I31({right_width_0_height_1_subtile_0__pin_I31_0_, right_width_0_height_1_subtile_0__pin_I31_1_, right_width_0_height_1_subtile_0__pin_I31_2_, right_width_0_height_1_subtile_0__pin_I31_3_, right_width_0_height_1_subtile_0__pin_I31_4_, right_width_0_height_1_subtile_0__pin_I31_5_, right_width_0_height_1_subtile_0__pin_I31_6_, right_width_0_height_1_subtile_0__pin_I31_7_, right_width_0_height_1_subtile_0__pin_I31_8_, right_width_0_height_1_subtile_0__pin_I31_9_, right_width_0_height_1_subtile_0__pin_I31_10_, right_width_0_height_1_subtile_0__pin_I31_11_}),
		.bram_IS1({top_width_0_height_1_subtile_0__pin_IS1_0_, top_width_0_height_1_subtile_0__pin_IS1_1_, top_width_0_height_1_subtile_0__pin_IS1_2_, right_width_0_height_1_subtile_0__pin_IS1_3_, right_width_0_height_1_subtile_0__pin_IS1_4_, right_width_0_height_1_subtile_0__pin_IS1_5_}),
		.bram_I02({top_width_0_height_2_subtile_0__pin_I02_0_, top_width_0_height_2_subtile_0__pin_I02_1_, top_width_0_height_2_subtile_0__pin_I02_2_, top_width_0_height_2_subtile_0__pin_I02_3_, top_width_0_height_2_subtile_0__pin_I02_4_, top_width_0_height_2_subtile_0__pin_I02_5_, top_width_0_height_2_subtile_0__pin_I02_6_, top_width_0_height_2_subtile_0__pin_I02_7_, top_width_0_height_2_subtile_0__pin_I02_8_, top_width_0_height_2_subtile_0__pin_I02_9_, top_width_0_height_2_subtile_0__pin_I02_10_, top_width_0_height_2_subtile_0__pin_I02_11_}),
		.bram_I12({top_width_0_height_2_subtile_0__pin_I12_0_, top_width_0_height_2_subtile_0__pin_I12_1_, top_width_0_height_2_subtile_0__pin_I12_2_, top_width_0_height_2_subtile_0__pin_I12_3_, top_width_0_height_2_subtile_0__pin_I12_4_, top_width_0_height_2_subtile_0__pin_I12_5_, top_width_0_height_2_subtile_0__pin_I12_6_, top_width_0_height_2_subtile_0__pin_I12_7_, top_width_0_height_2_subtile_0__pin_I12_8_, top_width_0_height_2_subtile_0__pin_I12_9_, top_width_0_height_2_subtile_0__pin_I12_10_, top_width_0_height_2_subtile_0__pin_I12_11_}),
		.bram_I22({right_width_0_height_2_subtile_0__pin_I22_0_, right_width_0_height_2_subtile_0__pin_I22_1_, right_width_0_height_2_subtile_0__pin_I22_2_, right_width_0_height_2_subtile_0__pin_I22_3_, right_width_0_height_2_subtile_0__pin_I22_4_, right_width_0_height_2_subtile_0__pin_I22_5_, right_width_0_height_2_subtile_0__pin_I22_6_, right_width_0_height_2_subtile_0__pin_I22_7_, right_width_0_height_2_subtile_0__pin_I22_8_, right_width_0_height_2_subtile_0__pin_I22_9_, right_width_0_height_2_subtile_0__pin_I22_10_, right_width_0_height_2_subtile_0__pin_I22_11_}),
		.bram_I32({right_width_0_height_2_subtile_0__pin_I32_0_, right_width_0_height_2_subtile_0__pin_I32_1_, right_width_0_height_2_subtile_0__pin_I32_2_, right_width_0_height_2_subtile_0__pin_I32_3_, right_width_0_height_2_subtile_0__pin_I32_4_, right_width_0_height_2_subtile_0__pin_I32_5_, right_width_0_height_2_subtile_0__pin_I32_6_, right_width_0_height_2_subtile_0__pin_I32_7_, right_width_0_height_2_subtile_0__pin_I32_8_, right_width_0_height_2_subtile_0__pin_I32_9_, right_width_0_height_2_subtile_0__pin_I32_10_, right_width_0_height_2_subtile_0__pin_I32_11_}),
		.bram_IS2({top_width_0_height_2_subtile_0__pin_IS2_0_, top_width_0_height_2_subtile_0__pin_IS2_1_, top_width_0_height_2_subtile_0__pin_IS2_2_, right_width_0_height_2_subtile_0__pin_IS2_3_, right_width_0_height_2_subtile_0__pin_IS2_4_, right_width_0_height_2_subtile_0__pin_IS2_5_}),
		.bram_sc_in({left_width_0_height_0_subtile_0__pin_sc_in_0_, left_width_0_height_0_subtile_0__pin_sc_in_1_, left_width_0_height_0_subtile_0__pin_sc_in_2_, left_width_0_height_0_subtile_0__pin_sc_in_3_, left_width_0_height_0_subtile_0__pin_sc_in_4_, left_width_0_height_0_subtile_0__pin_sc_in_5_, left_width_0_height_0_subtile_0__pin_sc_in_6_, left_width_0_height_0_subtile_0__pin_sc_in_7_, left_width_0_height_0_subtile_0__pin_sc_in_8_, left_width_0_height_0_subtile_0__pin_sc_in_9_, left_width_0_height_0_subtile_0__pin_sc_in_10_, left_width_0_height_0_subtile_0__pin_sc_in_11_, left_width_0_height_0_subtile_0__pin_sc_in_12_, left_width_0_height_0_subtile_0__pin_sc_in_13_, left_width_0_height_0_subtile_0__pin_sc_in_14_, left_width_0_height_0_subtile_0__pin_sc_in_15_, left_width_0_height_0_subtile_0__pin_sc_in_16_, left_width_0_height_0_subtile_0__pin_sc_in_17_, left_width_0_height_0_subtile_0__pin_sc_in_18_, left_width_0_height_0_subtile_0__pin_sc_in_19_, left_width_0_height_0_subtile_0__pin_sc_in_20_, left_width_0_height_0_subtile_0__pin_sc_in_21_, left_width_0_height_0_subtile_0__pin_sc_in_22_, left_width_0_height_0_subtile_0__pin_sc_in_23_, left_width_0_height_0_subtile_0__pin_sc_in_24_, left_width_0_height_0_subtile_0__pin_sc_in_25_, left_width_0_height_0_subtile_0__pin_sc_in_26_, left_width_0_height_0_subtile_0__pin_sc_in_27_, left_width_0_height_0_subtile_0__pin_sc_in_28_, left_width_0_height_0_subtile_0__pin_sc_in_29_, left_width_0_height_0_subtile_0__pin_sc_in_30_, left_width_0_height_0_subtile_0__pin_sc_in_31_, left_width_0_height_0_subtile_0__pin_sc_in_32_, left_width_0_height_0_subtile_0__pin_sc_in_33_, left_width_0_height_0_subtile_0__pin_sc_in_34_, left_width_0_height_0_subtile_0__pin_sc_in_35_, left_width_0_height_0_subtile_0__pin_sc_in_36_, left_width_0_height_0_subtile_0__pin_sc_in_37_, left_width_0_height_0_subtile_0__pin_sc_in_38_, left_width_0_height_0_subtile_0__pin_sc_in_39_, left_width_0_height_0_subtile_0__pin_sc_in_40_, left_width_0_height_0_subtile_0__pin_sc_in_41_, left_width_0_height_0_subtile_0__pin_sc_in_42_, left_width_0_height_0_subtile_0__pin_sc_in_43_, left_width_0_height_0_subtile_0__pin_sc_in_44_, left_width_0_height_0_subtile_0__pin_sc_in_45_, left_width_0_height_0_subtile_0__pin_sc_in_46_, left_width_0_height_0_subtile_0__pin_sc_in_47_}),
		.bram_RAM_ID_i({left_width_0_height_1_subtile_0__pin_RAM_ID_i_0_, left_width_0_height_1_subtile_0__pin_RAM_ID_i_1_, left_width_0_height_1_subtile_0__pin_RAM_ID_i_2_, left_width_0_height_1_subtile_0__pin_RAM_ID_i_3_, left_width_0_height_1_subtile_0__pin_RAM_ID_i_4_, left_width_0_height_1_subtile_0__pin_RAM_ID_i_5_, left_width_0_height_1_subtile_0__pin_RAM_ID_i_6_, left_width_0_height_1_subtile_0__pin_RAM_ID_i_7_, left_width_0_height_1_subtile_0__pin_RAM_ID_i_8_, left_width_0_height_1_subtile_0__pin_RAM_ID_i_9_, left_width_0_height_1_subtile_0__pin_RAM_ID_i_10_, left_width_0_height_1_subtile_0__pin_RAM_ID_i_11_, left_width_0_height_1_subtile_0__pin_RAM_ID_i_12_, left_width_0_height_1_subtile_0__pin_RAM_ID_i_13_, left_width_0_height_1_subtile_0__pin_RAM_ID_i_14_, left_width_0_height_1_subtile_0__pin_RAM_ID_i_15_, left_width_0_height_1_subtile_0__pin_RAM_ID_i_16_, left_width_0_height_1_subtile_0__pin_RAM_ID_i_17_, left_width_0_height_1_subtile_0__pin_RAM_ID_i_18_, left_width_0_height_1_subtile_0__pin_RAM_ID_i_19_}),
		.bram_PL_IN({top_width_0_height_2_subtile_0__pin_PL_IN_0_, top_width_0_height_2_subtile_0__pin_PL_IN_1_, top_width_0_height_2_subtile_0__pin_PL_IN_2_, top_width_0_height_2_subtile_0__pin_PL_IN_3_, top_width_0_height_2_subtile_0__pin_PL_IN_4_, top_width_0_height_2_subtile_0__pin_PL_IN_5_, top_width_0_height_2_subtile_0__pin_PL_IN_6_, top_width_0_height_2_subtile_0__pin_PL_IN_7_, top_width_0_height_2_subtile_0__pin_PL_IN_8_, top_width_0_height_2_subtile_0__pin_PL_IN_9_, top_width_0_height_2_subtile_0__pin_PL_IN_10_, top_width_0_height_2_subtile_0__pin_PL_IN_11_, top_width_0_height_2_subtile_0__pin_PL_IN_12_, top_width_0_height_2_subtile_0__pin_PL_IN_13_, top_width_0_height_2_subtile_0__pin_PL_IN_14_, top_width_0_height_2_subtile_0__pin_PL_IN_15_, top_width_0_height_2_subtile_0__pin_PL_IN_16_, top_width_0_height_2_subtile_0__pin_PL_IN_17_, top_width_0_height_2_subtile_0__pin_PL_IN_18_, top_width_0_height_2_subtile_0__pin_PL_IN_19_, top_width_0_height_2_subtile_0__pin_PL_IN_20_, top_width_0_height_2_subtile_0__pin_PL_IN_21_, top_width_0_height_2_subtile_0__pin_PL_IN_22_, top_width_0_height_2_subtile_0__pin_PL_IN_23_, top_width_0_height_2_subtile_0__pin_PL_IN_24_, top_width_0_height_2_subtile_0__pin_PL_IN_25_, top_width_0_height_2_subtile_0__pin_PL_IN_26_, top_width_0_height_2_subtile_0__pin_PL_IN_27_, top_width_0_height_2_subtile_0__pin_PL_IN_28_, top_width_0_height_2_subtile_0__pin_PL_IN_29_, top_width_0_height_2_subtile_0__pin_PL_IN_30_, top_width_0_height_2_subtile_0__pin_PL_IN_31_, top_width_0_height_2_subtile_0__pin_PL_IN_32_, top_width_0_height_2_subtile_0__pin_PL_IN_33_, top_width_0_height_2_subtile_0__pin_PL_IN_34_, top_width_0_height_2_subtile_0__pin_PL_IN_35_, top_width_0_height_2_subtile_0__pin_PL_IN_36_, top_width_0_height_2_subtile_0__pin_PL_IN_37_, top_width_0_height_2_subtile_0__pin_PL_IN_38_, top_width_0_height_2_subtile_0__pin_PL_IN_39_, top_width_0_height_2_subtile_0__pin_PL_IN_40_, top_width_0_height_2_subtile_0__pin_PL_IN_41_, top_width_0_height_2_subtile_0__pin_PL_IN_42_, top_width_0_height_2_subtile_0__pin_PL_IN_43_, top_width_0_height_2_subtile_0__pin_PL_IN_44_, top_width_0_height_2_subtile_0__pin_PL_IN_45_, top_width_0_height_2_subtile_0__pin_PL_IN_46_, top_width_0_height_2_subtile_0__pin_PL_IN_47_, top_width_0_height_2_subtile_0__pin_PL_IN_48_, top_width_0_height_2_subtile_0__pin_PL_IN_49_, top_width_0_height_2_subtile_0__pin_PL_IN_50_, top_width_0_height_2_subtile_0__pin_PL_IN_51_, top_width_0_height_2_subtile_0__pin_PL_IN_52_, top_width_0_height_2_subtile_0__pin_PL_IN_53_, top_width_0_height_2_subtile_0__pin_PL_IN_54_, top_width_0_height_2_subtile_0__pin_PL_IN_55_, top_width_0_height_2_subtile_0__pin_PL_IN_56_, top_width_0_height_2_subtile_0__pin_PL_IN_57_, top_width_0_height_2_subtile_0__pin_PL_IN_58_, top_width_0_height_2_subtile_0__pin_PL_IN_59_, top_width_0_height_2_subtile_0__pin_PL_IN_60_, top_width_0_height_2_subtile_0__pin_PL_IN_61_, top_width_0_height_2_subtile_0__pin_PL_IN_62_, top_width_0_height_2_subtile_0__pin_PL_IN_63_, top_width_0_height_2_subtile_0__pin_PL_IN_64_, top_width_0_height_2_subtile_0__pin_PL_IN_65_, top_width_0_height_2_subtile_0__pin_PL_IN_66_, top_width_0_height_2_subtile_0__pin_PL_IN_67_, top_width_0_height_2_subtile_0__pin_PL_IN_68_, top_width_0_height_2_subtile_0__pin_PL_IN_69_, top_width_0_height_2_subtile_0__pin_PL_IN_70_, top_width_0_height_2_subtile_0__pin_PL_IN_71_, top_width_0_height_2_subtile_0__pin_PL_IN_72_, top_width_0_height_2_subtile_0__pin_PL_IN_73_}),
		.bram_PL_DATA_IN({bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_0_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_1_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_2_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_3_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_4_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_5_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_6_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_7_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_8_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_9_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_10_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_11_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_12_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_13_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_14_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_15_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_16_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_17_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_18_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_19_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_20_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_21_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_22_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_23_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_24_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_25_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_26_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_27_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_28_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_29_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_30_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_31_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_32_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_33_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_34_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_IN_35_}),
		.bram_clk({left_width_0_height_0_subtile_0__pin_clk_0_, left_width_0_height_0_subtile_0__pin_clk_1_, left_width_0_height_0_subtile_0__pin_clk_2_, left_width_0_height_0_subtile_0__pin_clk_3_, left_width_0_height_0_subtile_0__pin_clk_4_, left_width_0_height_0_subtile_0__pin_clk_5_, left_width_0_height_0_subtile_0__pin_clk_6_, left_width_0_height_0_subtile_0__pin_clk_7_, left_width_0_height_0_subtile_0__pin_clk_8_, left_width_0_height_0_subtile_0__pin_clk_9_, left_width_0_height_0_subtile_0__pin_clk_10_, left_width_0_height_0_subtile_0__pin_clk_11_, left_width_0_height_0_subtile_0__pin_clk_12_, left_width_0_height_0_subtile_0__pin_clk_13_, left_width_0_height_0_subtile_0__pin_clk_14_, left_width_0_height_0_subtile_0__pin_clk_15_}),
		.ccff_head(ccff_head),
		.bram_O0({top_width_0_height_0_subtile_0__pin_O0_0_, top_width_0_height_0_subtile_0__pin_O0_1_, top_width_0_height_0_subtile_0__pin_O0_2_, top_width_0_height_0_subtile_0__pin_O0_3_, top_width_0_height_0_subtile_0__pin_O0_4_, top_width_0_height_0_subtile_0__pin_O0_5_, top_width_0_height_0_subtile_0__pin_O0_6_, top_width_0_height_0_subtile_0__pin_O0_7_, top_width_0_height_0_subtile_0__pin_O0_8_, top_width_0_height_0_subtile_0__pin_O0_9_, top_width_0_height_0_subtile_0__pin_O0_10_, top_width_0_height_0_subtile_0__pin_O0_11_, right_width_0_height_0_subtile_0__pin_O0_12_, right_width_0_height_0_subtile_0__pin_O0_13_, right_width_0_height_0_subtile_0__pin_O0_14_, right_width_0_height_0_subtile_0__pin_O0_15_, right_width_0_height_0_subtile_0__pin_O0_16_, right_width_0_height_0_subtile_0__pin_O0_17_, right_width_0_height_0_subtile_0__pin_O0_18_, right_width_0_height_0_subtile_0__pin_O0_19_, right_width_0_height_0_subtile_0__pin_O0_20_, right_width_0_height_0_subtile_0__pin_O0_21_, right_width_0_height_0_subtile_0__pin_O0_22_, right_width_0_height_0_subtile_0__pin_O0_23_}),
		.bram_O1({top_width_0_height_1_subtile_0__pin_O1_0_, top_width_0_height_1_subtile_0__pin_O1_1_, top_width_0_height_1_subtile_0__pin_O1_2_, top_width_0_height_1_subtile_0__pin_O1_3_, top_width_0_height_1_subtile_0__pin_O1_4_, top_width_0_height_1_subtile_0__pin_O1_5_, top_width_0_height_1_subtile_0__pin_O1_6_, top_width_0_height_1_subtile_0__pin_O1_7_, top_width_0_height_1_subtile_0__pin_O1_8_, top_width_0_height_1_subtile_0__pin_O1_9_, top_width_0_height_1_subtile_0__pin_O1_10_, top_width_0_height_1_subtile_0__pin_O1_11_, right_width_0_height_1_subtile_0__pin_O1_12_, right_width_0_height_1_subtile_0__pin_O1_13_, right_width_0_height_1_subtile_0__pin_O1_14_, right_width_0_height_1_subtile_0__pin_O1_15_, right_width_0_height_1_subtile_0__pin_O1_16_, right_width_0_height_1_subtile_0__pin_O1_17_, right_width_0_height_1_subtile_0__pin_O1_18_, right_width_0_height_1_subtile_0__pin_O1_19_, right_width_0_height_1_subtile_0__pin_O1_20_, right_width_0_height_1_subtile_0__pin_O1_21_, right_width_0_height_1_subtile_0__pin_O1_22_, right_width_0_height_1_subtile_0__pin_O1_23_}),
		.bram_O2({top_width_0_height_2_subtile_0__pin_O2_0_, top_width_0_height_2_subtile_0__pin_O2_1_, top_width_0_height_2_subtile_0__pin_O2_2_, top_width_0_height_2_subtile_0__pin_O2_3_, top_width_0_height_2_subtile_0__pin_O2_4_, top_width_0_height_2_subtile_0__pin_O2_5_, top_width_0_height_2_subtile_0__pin_O2_6_, top_width_0_height_2_subtile_0__pin_O2_7_, top_width_0_height_2_subtile_0__pin_O2_8_, top_width_0_height_2_subtile_0__pin_O2_9_, top_width_0_height_2_subtile_0__pin_O2_10_, top_width_0_height_2_subtile_0__pin_O2_11_, right_width_0_height_2_subtile_0__pin_O2_12_, right_width_0_height_2_subtile_0__pin_O2_13_, right_width_0_height_2_subtile_0__pin_O2_14_, right_width_0_height_2_subtile_0__pin_O2_15_, right_width_0_height_2_subtile_0__pin_O2_16_, right_width_0_height_2_subtile_0__pin_O2_17_, right_width_0_height_2_subtile_0__pin_O2_18_, right_width_0_height_2_subtile_0__pin_O2_19_, right_width_0_height_2_subtile_0__pin_O2_20_, right_width_0_height_2_subtile_0__pin_O2_21_, right_width_0_height_2_subtile_0__pin_O2_22_, right_width_0_height_2_subtile_0__pin_O2_23_}),
		.bram_sc_out({right_width_0_height_0_subtile_0__pin_sc_out_0_, right_width_0_height_0_subtile_0__pin_sc_out_1_, right_width_0_height_0_subtile_0__pin_sc_out_2_, right_width_0_height_0_subtile_0__pin_sc_out_3_, right_width_0_height_0_subtile_0__pin_sc_out_4_, right_width_0_height_0_subtile_0__pin_sc_out_5_, right_width_0_height_0_subtile_0__pin_sc_out_6_, right_width_0_height_0_subtile_0__pin_sc_out_7_, right_width_0_height_0_subtile_0__pin_sc_out_8_, right_width_0_height_0_subtile_0__pin_sc_out_9_, right_width_0_height_0_subtile_0__pin_sc_out_10_, right_width_0_height_0_subtile_0__pin_sc_out_11_, right_width_0_height_0_subtile_0__pin_sc_out_12_, right_width_0_height_0_subtile_0__pin_sc_out_13_, right_width_0_height_0_subtile_0__pin_sc_out_14_, right_width_0_height_0_subtile_0__pin_sc_out_15_, right_width_0_height_0_subtile_0__pin_sc_out_16_, right_width_0_height_0_subtile_0__pin_sc_out_17_, right_width_0_height_0_subtile_0__pin_sc_out_18_, right_width_0_height_0_subtile_0__pin_sc_out_19_, right_width_0_height_0_subtile_0__pin_sc_out_20_, right_width_0_height_0_subtile_0__pin_sc_out_21_, right_width_0_height_0_subtile_0__pin_sc_out_22_, right_width_0_height_0_subtile_0__pin_sc_out_23_, right_width_0_height_0_subtile_0__pin_sc_out_24_, right_width_0_height_0_subtile_0__pin_sc_out_25_, right_width_0_height_0_subtile_0__pin_sc_out_26_, right_width_0_height_0_subtile_0__pin_sc_out_27_, right_width_0_height_0_subtile_0__pin_sc_out_28_, right_width_0_height_0_subtile_0__pin_sc_out_29_, right_width_0_height_0_subtile_0__pin_sc_out_30_, right_width_0_height_0_subtile_0__pin_sc_out_31_, right_width_0_height_0_subtile_0__pin_sc_out_32_, right_width_0_height_0_subtile_0__pin_sc_out_33_, right_width_0_height_0_subtile_0__pin_sc_out_34_, right_width_0_height_0_subtile_0__pin_sc_out_35_, right_width_0_height_0_subtile_0__pin_sc_out_36_, right_width_0_height_0_subtile_0__pin_sc_out_37_, right_width_0_height_0_subtile_0__pin_sc_out_38_, right_width_0_height_0_subtile_0__pin_sc_out_39_, right_width_0_height_0_subtile_0__pin_sc_out_40_, right_width_0_height_0_subtile_0__pin_sc_out_41_, right_width_0_height_0_subtile_0__pin_sc_out_42_, right_width_0_height_0_subtile_0__pin_sc_out_43_, right_width_0_height_0_subtile_0__pin_sc_out_44_, right_width_0_height_0_subtile_0__pin_sc_out_45_, right_width_0_height_0_subtile_0__pin_sc_out_46_, right_width_0_height_0_subtile_0__pin_sc_out_47_}),
		.bram_PL_OUT({bottom_width_0_height_0_subtile_0__pin_PL_OUT_0_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_1_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_2_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_3_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_4_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_5_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_6_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_7_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_8_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_9_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_10_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_11_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_12_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_13_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_14_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_15_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_16_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_17_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_18_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_19_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_20_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_21_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_22_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_23_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_24_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_25_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_26_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_27_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_28_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_29_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_30_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_31_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_32_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_33_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_34_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_35_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_36_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_37_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_38_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_39_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_40_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_41_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_42_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_43_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_44_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_45_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_46_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_47_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_48_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_49_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_50_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_51_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_52_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_53_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_54_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_55_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_56_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_57_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_58_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_59_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_60_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_61_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_62_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_63_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_64_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_65_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_66_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_67_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_68_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_69_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_70_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_71_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_72_, bottom_width_0_height_0_subtile_0__pin_PL_OUT_73_}),
		.bram_PL_DATA_OUT({top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_0_, top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_1_, top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_2_, top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_3_, top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_4_, top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_5_, top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_6_, top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_7_, top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_8_, top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_9_, top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_10_, top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_11_, top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_12_, top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_13_, top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_14_, top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_15_, top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_16_, top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_17_, top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_18_, top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_19_, top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_20_, top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_21_, top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_22_, top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_23_, top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_24_, top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_25_, top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_26_, top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_27_, top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_28_, top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_29_, top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_30_, top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_31_, top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_32_, top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_33_, top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_34_, top_width_0_height_2_subtile_0__pin_PL_DATA_OUT_35_}),
		.ccff_tail(ccff_tail));

endmodule
// ----- END Verilog module for grid_bram -----

//----- Default net type -----
`default_nettype none



// ----- END Grid Verilog module: grid_bram -----

