//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for physical tile: dsp]
//	Author: Xifan TANG
//	Organization: University of Utah
//-------------------------------------------
//----- Time scale -----
`timescale 1ns / 1ps

// ----- BEGIN Grid Verilog module: grid_dsp -----
//----- Default net type -----
`default_nettype wire

// ----- Verilog module for grid_dsp -----
module grid_dsp(scan_mode,
                scan_enable,
                global_reset,
                config_enable,
                prog_clock,
                top_width_0_height_0_subtile_0__pin_I00_0_,
                top_width_0_height_0_subtile_0__pin_I00_1_,
                top_width_0_height_0_subtile_0__pin_I00_2_,
                top_width_0_height_0_subtile_0__pin_I00_3_,
                top_width_0_height_0_subtile_0__pin_I00_4_,
                top_width_0_height_0_subtile_0__pin_I00_5_,
                top_width_0_height_0_subtile_0__pin_I00_6_,
                top_width_0_height_0_subtile_0__pin_I00_7_,
                top_width_0_height_0_subtile_0__pin_I00_8_,
                top_width_0_height_0_subtile_0__pin_I00_9_,
                top_width_0_height_0_subtile_0__pin_I00_10_,
                top_width_0_height_0_subtile_0__pin_I00_11_,
                top_width_0_height_0_subtile_0__pin_I10_0_,
                top_width_0_height_0_subtile_0__pin_I10_1_,
                top_width_0_height_0_subtile_0__pin_I10_2_,
                top_width_0_height_0_subtile_0__pin_I10_3_,
                top_width_0_height_0_subtile_0__pin_I10_4_,
                top_width_0_height_0_subtile_0__pin_I10_5_,
                top_width_0_height_0_subtile_0__pin_I10_6_,
                top_width_0_height_0_subtile_0__pin_I10_7_,
                top_width_0_height_0_subtile_0__pin_I10_8_,
                top_width_0_height_0_subtile_0__pin_I10_9_,
                top_width_0_height_0_subtile_0__pin_I10_10_,
                top_width_0_height_0_subtile_0__pin_I10_11_,
                top_width_0_height_0_subtile_0__pin_IS0_0_,
                top_width_0_height_0_subtile_0__pin_IS0_1_,
                top_width_0_height_0_subtile_0__pin_IS0_2_,
                top_width_0_height_1_subtile_0__pin_I01_0_,
                top_width_0_height_1_subtile_0__pin_I01_1_,
                top_width_0_height_1_subtile_0__pin_I01_2_,
                top_width_0_height_1_subtile_0__pin_I01_3_,
                top_width_0_height_1_subtile_0__pin_I01_4_,
                top_width_0_height_1_subtile_0__pin_I01_5_,
                top_width_0_height_1_subtile_0__pin_I01_6_,
                top_width_0_height_1_subtile_0__pin_I01_7_,
                top_width_0_height_1_subtile_0__pin_I01_8_,
                top_width_0_height_1_subtile_0__pin_I01_9_,
                top_width_0_height_1_subtile_0__pin_I01_10_,
                top_width_0_height_1_subtile_0__pin_I01_11_,
                top_width_0_height_1_subtile_0__pin_I11_0_,
                top_width_0_height_1_subtile_0__pin_I11_1_,
                top_width_0_height_1_subtile_0__pin_I11_2_,
                top_width_0_height_1_subtile_0__pin_I11_3_,
                top_width_0_height_1_subtile_0__pin_I11_4_,
                top_width_0_height_1_subtile_0__pin_I11_5_,
                top_width_0_height_1_subtile_0__pin_I11_6_,
                top_width_0_height_1_subtile_0__pin_I11_7_,
                top_width_0_height_1_subtile_0__pin_I11_8_,
                top_width_0_height_1_subtile_0__pin_I11_9_,
                top_width_0_height_1_subtile_0__pin_I11_10_,
                top_width_0_height_1_subtile_0__pin_I11_11_,
                top_width_0_height_1_subtile_0__pin_IS1_0_,
                top_width_0_height_1_subtile_0__pin_IS1_1_,
                top_width_0_height_1_subtile_0__pin_IS1_2_,
                top_width_0_height_2_subtile_0__pin_I02_0_,
                top_width_0_height_2_subtile_0__pin_I02_1_,
                top_width_0_height_2_subtile_0__pin_I02_2_,
                top_width_0_height_2_subtile_0__pin_I02_3_,
                top_width_0_height_2_subtile_0__pin_I02_4_,
                top_width_0_height_2_subtile_0__pin_I02_5_,
                top_width_0_height_2_subtile_0__pin_I02_6_,
                top_width_0_height_2_subtile_0__pin_I02_7_,
                top_width_0_height_2_subtile_0__pin_I02_8_,
                top_width_0_height_2_subtile_0__pin_I02_9_,
                top_width_0_height_2_subtile_0__pin_I02_10_,
                top_width_0_height_2_subtile_0__pin_I02_11_,
                top_width_0_height_2_subtile_0__pin_I12_0_,
                top_width_0_height_2_subtile_0__pin_I12_1_,
                top_width_0_height_2_subtile_0__pin_I12_2_,
                top_width_0_height_2_subtile_0__pin_I12_3_,
                top_width_0_height_2_subtile_0__pin_I12_4_,
                top_width_0_height_2_subtile_0__pin_I12_5_,
                top_width_0_height_2_subtile_0__pin_I12_6_,
                top_width_0_height_2_subtile_0__pin_I12_7_,
                top_width_0_height_2_subtile_0__pin_I12_8_,
                top_width_0_height_2_subtile_0__pin_I12_9_,
                top_width_0_height_2_subtile_0__pin_I12_10_,
                top_width_0_height_2_subtile_0__pin_I12_11_,
                top_width_0_height_2_subtile_0__pin_IS2_0_,
                top_width_0_height_2_subtile_0__pin_IS2_1_,
                top_width_0_height_2_subtile_0__pin_IS2_2_,
                right_width_0_height_0_subtile_0__pin_I20_0_,
                right_width_0_height_0_subtile_0__pin_I20_1_,
                right_width_0_height_0_subtile_0__pin_I20_2_,
                right_width_0_height_0_subtile_0__pin_I20_3_,
                right_width_0_height_0_subtile_0__pin_I20_4_,
                right_width_0_height_0_subtile_0__pin_I20_5_,
                right_width_0_height_0_subtile_0__pin_I20_6_,
                right_width_0_height_0_subtile_0__pin_I20_7_,
                right_width_0_height_0_subtile_0__pin_I20_8_,
                right_width_0_height_0_subtile_0__pin_I20_9_,
                right_width_0_height_0_subtile_0__pin_I20_10_,
                right_width_0_height_0_subtile_0__pin_I20_11_,
                right_width_0_height_0_subtile_0__pin_I30_0_,
                right_width_0_height_0_subtile_0__pin_I30_1_,
                right_width_0_height_0_subtile_0__pin_I30_2_,
                right_width_0_height_0_subtile_0__pin_I30_3_,
                right_width_0_height_0_subtile_0__pin_I30_4_,
                right_width_0_height_0_subtile_0__pin_I30_5_,
                right_width_0_height_0_subtile_0__pin_I30_6_,
                right_width_0_height_0_subtile_0__pin_I30_7_,
                right_width_0_height_0_subtile_0__pin_I30_8_,
                right_width_0_height_0_subtile_0__pin_I30_9_,
                right_width_0_height_0_subtile_0__pin_I30_10_,
                right_width_0_height_0_subtile_0__pin_I30_11_,
                right_width_0_height_0_subtile_0__pin_IS0_3_,
                right_width_0_height_0_subtile_0__pin_IS0_4_,
                right_width_0_height_0_subtile_0__pin_IS0_5_,
                right_width_0_height_1_subtile_0__pin_I21_0_,
                right_width_0_height_1_subtile_0__pin_I21_1_,
                right_width_0_height_1_subtile_0__pin_I21_2_,
                right_width_0_height_1_subtile_0__pin_I21_3_,
                right_width_0_height_1_subtile_0__pin_I21_4_,
                right_width_0_height_1_subtile_0__pin_I21_5_,
                right_width_0_height_1_subtile_0__pin_I21_6_,
                right_width_0_height_1_subtile_0__pin_I21_7_,
                right_width_0_height_1_subtile_0__pin_I21_8_,
                right_width_0_height_1_subtile_0__pin_I21_9_,
                right_width_0_height_1_subtile_0__pin_I21_10_,
                right_width_0_height_1_subtile_0__pin_I21_11_,
                right_width_0_height_1_subtile_0__pin_I31_0_,
                right_width_0_height_1_subtile_0__pin_I31_1_,
                right_width_0_height_1_subtile_0__pin_I31_2_,
                right_width_0_height_1_subtile_0__pin_I31_3_,
                right_width_0_height_1_subtile_0__pin_I31_4_,
                right_width_0_height_1_subtile_0__pin_I31_5_,
                right_width_0_height_1_subtile_0__pin_I31_6_,
                right_width_0_height_1_subtile_0__pin_I31_7_,
                right_width_0_height_1_subtile_0__pin_I31_8_,
                right_width_0_height_1_subtile_0__pin_I31_9_,
                right_width_0_height_1_subtile_0__pin_I31_10_,
                right_width_0_height_1_subtile_0__pin_I31_11_,
                right_width_0_height_1_subtile_0__pin_IS1_3_,
                right_width_0_height_1_subtile_0__pin_IS1_4_,
                right_width_0_height_1_subtile_0__pin_IS1_5_,
                right_width_0_height_2_subtile_0__pin_I22_0_,
                right_width_0_height_2_subtile_0__pin_I22_1_,
                right_width_0_height_2_subtile_0__pin_I22_2_,
                right_width_0_height_2_subtile_0__pin_I22_3_,
                right_width_0_height_2_subtile_0__pin_I22_4_,
                right_width_0_height_2_subtile_0__pin_I22_5_,
                right_width_0_height_2_subtile_0__pin_I22_6_,
                right_width_0_height_2_subtile_0__pin_I22_7_,
                right_width_0_height_2_subtile_0__pin_I22_8_,
                right_width_0_height_2_subtile_0__pin_I22_9_,
                right_width_0_height_2_subtile_0__pin_I22_10_,
                right_width_0_height_2_subtile_0__pin_I22_11_,
                right_width_0_height_2_subtile_0__pin_I32_0_,
                right_width_0_height_2_subtile_0__pin_I32_1_,
                right_width_0_height_2_subtile_0__pin_I32_2_,
                right_width_0_height_2_subtile_0__pin_I32_3_,
                right_width_0_height_2_subtile_0__pin_I32_4_,
                right_width_0_height_2_subtile_0__pin_I32_5_,
                right_width_0_height_2_subtile_0__pin_I32_6_,
                right_width_0_height_2_subtile_0__pin_I32_7_,
                right_width_0_height_2_subtile_0__pin_I32_8_,
                right_width_0_height_2_subtile_0__pin_I32_9_,
                right_width_0_height_2_subtile_0__pin_I32_10_,
                right_width_0_height_2_subtile_0__pin_I32_11_,
                right_width_0_height_2_subtile_0__pin_IS2_3_,
                right_width_0_height_2_subtile_0__pin_IS2_4_,
                right_width_0_height_2_subtile_0__pin_IS2_5_,
                left_width_0_height_0_subtile_0__pin_sc_in_0_,
                left_width_0_height_0_subtile_0__pin_sc_in_1_,
                left_width_0_height_0_subtile_0__pin_sc_in_2_,
                left_width_0_height_0_subtile_0__pin_sc_in_3_,
                left_width_0_height_0_subtile_0__pin_sc_in_4_,
                left_width_0_height_0_subtile_0__pin_sc_in_5_,
                left_width_0_height_0_subtile_0__pin_sc_in_6_,
                left_width_0_height_0_subtile_0__pin_sc_in_7_,
                left_width_0_height_0_subtile_0__pin_sc_in_8_,
                left_width_0_height_0_subtile_0__pin_sc_in_9_,
                left_width_0_height_0_subtile_0__pin_sc_in_10_,
                left_width_0_height_0_subtile_0__pin_sc_in_11_,
                left_width_0_height_0_subtile_0__pin_sc_in_12_,
                left_width_0_height_0_subtile_0__pin_sc_in_13_,
                left_width_0_height_0_subtile_0__pin_sc_in_14_,
                left_width_0_height_0_subtile_0__pin_sc_in_15_,
                left_width_0_height_0_subtile_0__pin_sc_in_16_,
                left_width_0_height_0_subtile_0__pin_sc_in_17_,
                left_width_0_height_0_subtile_0__pin_sc_in_18_,
                left_width_0_height_0_subtile_0__pin_sc_in_19_,
                left_width_0_height_0_subtile_0__pin_clk_0_,
                left_width_0_height_0_subtile_0__pin_clk_1_,
                left_width_0_height_0_subtile_0__pin_clk_2_,
                left_width_0_height_0_subtile_0__pin_clk_3_,
                left_width_0_height_0_subtile_0__pin_clk_4_,
                left_width_0_height_0_subtile_0__pin_clk_5_,
                left_width_0_height_0_subtile_0__pin_clk_6_,
                left_width_0_height_0_subtile_0__pin_clk_7_,
                left_width_0_height_0_subtile_0__pin_clk_8_,
                left_width_0_height_0_subtile_0__pin_clk_9_,
                left_width_0_height_0_subtile_0__pin_clk_10_,
                left_width_0_height_0_subtile_0__pin_clk_11_,
                left_width_0_height_0_subtile_0__pin_clk_12_,
                left_width_0_height_0_subtile_0__pin_clk_13_,
                left_width_0_height_0_subtile_0__pin_clk_14_,
                left_width_0_height_0_subtile_0__pin_clk_15_,
                ccff_head,
                top_width_0_height_0_subtile_0__pin_O0_0_,
                top_width_0_height_0_subtile_0__pin_O0_1_,
                top_width_0_height_0_subtile_0__pin_O0_2_,
                top_width_0_height_0_subtile_0__pin_O0_3_,
                top_width_0_height_0_subtile_0__pin_O0_4_,
                top_width_0_height_0_subtile_0__pin_O0_5_,
                top_width_0_height_0_subtile_0__pin_O0_6_,
                top_width_0_height_0_subtile_0__pin_O0_7_,
                top_width_0_height_0_subtile_0__pin_O0_8_,
                top_width_0_height_0_subtile_0__pin_O0_9_,
                top_width_0_height_0_subtile_0__pin_O0_10_,
                top_width_0_height_0_subtile_0__pin_O0_11_,
                top_width_0_height_1_subtile_0__pin_O1_0_,
                top_width_0_height_1_subtile_0__pin_O1_1_,
                top_width_0_height_1_subtile_0__pin_O1_2_,
                top_width_0_height_1_subtile_0__pin_O1_3_,
                top_width_0_height_1_subtile_0__pin_O1_4_,
                top_width_0_height_1_subtile_0__pin_O1_5_,
                top_width_0_height_1_subtile_0__pin_O1_6_,
                top_width_0_height_1_subtile_0__pin_O1_7_,
                top_width_0_height_1_subtile_0__pin_O1_8_,
                top_width_0_height_1_subtile_0__pin_O1_9_,
                top_width_0_height_1_subtile_0__pin_O1_10_,
                top_width_0_height_1_subtile_0__pin_O1_11_,
                top_width_0_height_2_subtile_0__pin_O2_0_,
                top_width_0_height_2_subtile_0__pin_O2_1_,
                top_width_0_height_2_subtile_0__pin_O2_2_,
                top_width_0_height_2_subtile_0__pin_O2_3_,
                top_width_0_height_2_subtile_0__pin_O2_4_,
                top_width_0_height_2_subtile_0__pin_O2_5_,
                top_width_0_height_2_subtile_0__pin_O2_6_,
                top_width_0_height_2_subtile_0__pin_O2_7_,
                top_width_0_height_2_subtile_0__pin_O2_8_,
                top_width_0_height_2_subtile_0__pin_O2_9_,
                top_width_0_height_2_subtile_0__pin_O2_10_,
                top_width_0_height_2_subtile_0__pin_O2_11_,
                right_width_0_height_0_subtile_0__pin_O0_12_,
                right_width_0_height_0_subtile_0__pin_O0_13_,
                right_width_0_height_0_subtile_0__pin_O0_14_,
                right_width_0_height_0_subtile_0__pin_O0_15_,
                right_width_0_height_0_subtile_0__pin_O0_16_,
                right_width_0_height_0_subtile_0__pin_O0_17_,
                right_width_0_height_0_subtile_0__pin_O0_18_,
                right_width_0_height_0_subtile_0__pin_O0_19_,
                right_width_0_height_0_subtile_0__pin_O0_20_,
                right_width_0_height_0_subtile_0__pin_O0_21_,
                right_width_0_height_0_subtile_0__pin_O0_22_,
                right_width_0_height_0_subtile_0__pin_O0_23_,
                right_width_0_height_0_subtile_0__pin_sc_out_0_,
                right_width_0_height_0_subtile_0__pin_sc_out_1_,
                right_width_0_height_0_subtile_0__pin_sc_out_2_,
                right_width_0_height_0_subtile_0__pin_sc_out_3_,
                right_width_0_height_0_subtile_0__pin_sc_out_4_,
                right_width_0_height_0_subtile_0__pin_sc_out_5_,
                right_width_0_height_0_subtile_0__pin_sc_out_6_,
                right_width_0_height_0_subtile_0__pin_sc_out_7_,
                right_width_0_height_0_subtile_0__pin_sc_out_8_,
                right_width_0_height_0_subtile_0__pin_sc_out_9_,
                right_width_0_height_0_subtile_0__pin_sc_out_10_,
                right_width_0_height_0_subtile_0__pin_sc_out_11_,
                right_width_0_height_0_subtile_0__pin_sc_out_12_,
                right_width_0_height_0_subtile_0__pin_sc_out_13_,
                right_width_0_height_0_subtile_0__pin_sc_out_14_,
                right_width_0_height_0_subtile_0__pin_sc_out_15_,
                right_width_0_height_0_subtile_0__pin_sc_out_16_,
                right_width_0_height_0_subtile_0__pin_sc_out_17_,
                right_width_0_height_0_subtile_0__pin_sc_out_18_,
                right_width_0_height_0_subtile_0__pin_sc_out_19_,
                right_width_0_height_1_subtile_0__pin_O1_12_,
                right_width_0_height_1_subtile_0__pin_O1_13_,
                right_width_0_height_1_subtile_0__pin_O1_14_,
                right_width_0_height_1_subtile_0__pin_O1_15_,
                right_width_0_height_1_subtile_0__pin_O1_16_,
                right_width_0_height_1_subtile_0__pin_O1_17_,
                right_width_0_height_1_subtile_0__pin_O1_18_,
                right_width_0_height_1_subtile_0__pin_O1_19_,
                right_width_0_height_1_subtile_0__pin_O1_20_,
                right_width_0_height_1_subtile_0__pin_O1_21_,
                right_width_0_height_1_subtile_0__pin_O1_22_,
                right_width_0_height_1_subtile_0__pin_O1_23_,
                right_width_0_height_2_subtile_0__pin_O2_12_,
                right_width_0_height_2_subtile_0__pin_O2_13_,
                right_width_0_height_2_subtile_0__pin_O2_14_,
                right_width_0_height_2_subtile_0__pin_O2_15_,
                right_width_0_height_2_subtile_0__pin_O2_16_,
                right_width_0_height_2_subtile_0__pin_O2_17_,
                right_width_0_height_2_subtile_0__pin_O2_18_,
                right_width_0_height_2_subtile_0__pin_O2_19_,
                right_width_0_height_2_subtile_0__pin_O2_20_,
                right_width_0_height_2_subtile_0__pin_O2_21_,
                right_width_0_height_2_subtile_0__pin_O2_22_,
                right_width_0_height_2_subtile_0__pin_O2_23_,
                ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] scan_mode;
//----- GLOBAL PORTS -----
input [0:0] scan_enable;
//----- GLOBAL PORTS -----
input [0:0] global_reset;
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_clock;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I00_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I00_1_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I00_2_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I00_3_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I00_4_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I00_5_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I00_6_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I00_7_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I00_8_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I00_9_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I00_10_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I00_11_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I10_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I10_1_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I10_2_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I10_3_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I10_4_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I10_5_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I10_6_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I10_7_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I10_8_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I10_9_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I10_10_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I10_11_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_IS0_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_IS0_1_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_IS0_2_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I01_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I01_1_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I01_2_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I01_3_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I01_4_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I01_5_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I01_6_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I01_7_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I01_8_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I01_9_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I01_10_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I01_11_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I11_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I11_1_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I11_2_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I11_3_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I11_4_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I11_5_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I11_6_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I11_7_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I11_8_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I11_9_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I11_10_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_I11_11_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_IS1_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_IS1_1_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_1_subtile_0__pin_IS1_2_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I02_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I02_1_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I02_2_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I02_3_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I02_4_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I02_5_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I02_6_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I02_7_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I02_8_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I02_9_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I02_10_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I02_11_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I12_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I12_1_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I12_2_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I12_3_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I12_4_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I12_5_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I12_6_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I12_7_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I12_8_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I12_9_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I12_10_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_I12_11_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_IS2_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_IS2_1_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_2_subtile_0__pin_IS2_2_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I20_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I20_1_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I20_2_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I20_3_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I20_4_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I20_5_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I20_6_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I20_7_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I20_8_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I20_9_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I20_10_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I20_11_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I30_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I30_1_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I30_2_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I30_3_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I30_4_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I30_5_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I30_6_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I30_7_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I30_8_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I30_9_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I30_10_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I30_11_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_IS0_3_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_IS0_4_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_IS0_5_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I21_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I21_1_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I21_2_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I21_3_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I21_4_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I21_5_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I21_6_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I21_7_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I21_8_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I21_9_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I21_10_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I21_11_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I31_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I31_1_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I31_2_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I31_3_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I31_4_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I31_5_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I31_6_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I31_7_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I31_8_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I31_9_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I31_10_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_I31_11_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_IS1_3_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_IS1_4_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_IS1_5_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I22_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I22_1_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I22_2_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I22_3_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I22_4_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I22_5_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I22_6_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I22_7_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I22_8_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I22_9_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I22_10_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I22_11_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I32_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I32_1_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I32_2_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I32_3_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I32_4_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I32_5_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I32_6_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I32_7_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I32_8_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I32_9_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I32_10_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_I32_11_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_IS2_3_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_IS2_4_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_IS2_5_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_1_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_2_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_3_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_4_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_5_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_6_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_7_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_8_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_9_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_10_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_11_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_12_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_13_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_14_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_15_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_16_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_17_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_18_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_19_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_O0_0_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_O0_1_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_O0_2_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_O0_3_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_O0_4_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_O0_5_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_O0_6_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_O0_7_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_O0_8_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_O0_9_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_O0_10_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_O0_11_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_1_subtile_0__pin_O1_0_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_1_subtile_0__pin_O1_1_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_1_subtile_0__pin_O1_2_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_1_subtile_0__pin_O1_3_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_1_subtile_0__pin_O1_4_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_1_subtile_0__pin_O1_5_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_1_subtile_0__pin_O1_6_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_1_subtile_0__pin_O1_7_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_1_subtile_0__pin_O1_8_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_1_subtile_0__pin_O1_9_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_1_subtile_0__pin_O1_10_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_1_subtile_0__pin_O1_11_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_O2_0_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_O2_1_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_O2_2_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_O2_3_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_O2_4_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_O2_5_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_O2_6_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_O2_7_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_O2_8_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_O2_9_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_O2_10_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_2_subtile_0__pin_O2_11_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_O0_12_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_O0_13_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_O0_14_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_O0_15_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_O0_16_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_O0_17_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_O0_18_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_O0_19_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_O0_20_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_O0_21_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_O0_22_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_O0_23_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_1_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_2_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_3_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_4_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_5_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_6_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_7_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_8_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_9_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_10_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_11_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_12_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_13_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_14_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_15_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_16_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_17_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_18_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_sc_out_19_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_O1_12_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_O1_13_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_O1_14_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_O1_15_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_O1_16_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_O1_17_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_O1_18_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_O1_19_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_O1_20_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_O1_21_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_O1_22_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_O1_23_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_2_subtile_0__pin_O2_12_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_2_subtile_0__pin_O2_13_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_2_subtile_0__pin_O2_14_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_2_subtile_0__pin_O2_15_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_2_subtile_0__pin_O2_16_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_2_subtile_0__pin_O2_17_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_2_subtile_0__pin_O2_18_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_2_subtile_0__pin_O2_19_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_2_subtile_0__pin_O2_20_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_2_subtile_0__pin_O2_21_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_2_subtile_0__pin_O2_22_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_2_subtile_0__pin_O2_23_;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	logical_tile_dsp_mode_dsp_ logical_tile_dsp_mode_dsp__0 (
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.global_reset(global_reset),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.dsp_I00({top_width_0_height_0_subtile_0__pin_I00_0_, top_width_0_height_0_subtile_0__pin_I00_1_, top_width_0_height_0_subtile_0__pin_I00_2_, top_width_0_height_0_subtile_0__pin_I00_3_, top_width_0_height_0_subtile_0__pin_I00_4_, top_width_0_height_0_subtile_0__pin_I00_5_, top_width_0_height_0_subtile_0__pin_I00_6_, top_width_0_height_0_subtile_0__pin_I00_7_, top_width_0_height_0_subtile_0__pin_I00_8_, top_width_0_height_0_subtile_0__pin_I00_9_, top_width_0_height_0_subtile_0__pin_I00_10_, top_width_0_height_0_subtile_0__pin_I00_11_}),
		.dsp_I10({top_width_0_height_0_subtile_0__pin_I10_0_, top_width_0_height_0_subtile_0__pin_I10_1_, top_width_0_height_0_subtile_0__pin_I10_2_, top_width_0_height_0_subtile_0__pin_I10_3_, top_width_0_height_0_subtile_0__pin_I10_4_, top_width_0_height_0_subtile_0__pin_I10_5_, top_width_0_height_0_subtile_0__pin_I10_6_, top_width_0_height_0_subtile_0__pin_I10_7_, top_width_0_height_0_subtile_0__pin_I10_8_, top_width_0_height_0_subtile_0__pin_I10_9_, top_width_0_height_0_subtile_0__pin_I10_10_, top_width_0_height_0_subtile_0__pin_I10_11_}),
		.dsp_I20({right_width_0_height_0_subtile_0__pin_I20_0_, right_width_0_height_0_subtile_0__pin_I20_1_, right_width_0_height_0_subtile_0__pin_I20_2_, right_width_0_height_0_subtile_0__pin_I20_3_, right_width_0_height_0_subtile_0__pin_I20_4_, right_width_0_height_0_subtile_0__pin_I20_5_, right_width_0_height_0_subtile_0__pin_I20_6_, right_width_0_height_0_subtile_0__pin_I20_7_, right_width_0_height_0_subtile_0__pin_I20_8_, right_width_0_height_0_subtile_0__pin_I20_9_, right_width_0_height_0_subtile_0__pin_I20_10_, right_width_0_height_0_subtile_0__pin_I20_11_}),
		.dsp_I30({right_width_0_height_0_subtile_0__pin_I30_0_, right_width_0_height_0_subtile_0__pin_I30_1_, right_width_0_height_0_subtile_0__pin_I30_2_, right_width_0_height_0_subtile_0__pin_I30_3_, right_width_0_height_0_subtile_0__pin_I30_4_, right_width_0_height_0_subtile_0__pin_I30_5_, right_width_0_height_0_subtile_0__pin_I30_6_, right_width_0_height_0_subtile_0__pin_I30_7_, right_width_0_height_0_subtile_0__pin_I30_8_, right_width_0_height_0_subtile_0__pin_I30_9_, right_width_0_height_0_subtile_0__pin_I30_10_, right_width_0_height_0_subtile_0__pin_I30_11_}),
		.dsp_IS0({top_width_0_height_0_subtile_0__pin_IS0_0_, top_width_0_height_0_subtile_0__pin_IS0_1_, top_width_0_height_0_subtile_0__pin_IS0_2_, right_width_0_height_0_subtile_0__pin_IS0_3_, right_width_0_height_0_subtile_0__pin_IS0_4_, right_width_0_height_0_subtile_0__pin_IS0_5_}),
		.dsp_I01({top_width_0_height_1_subtile_0__pin_I01_0_, top_width_0_height_1_subtile_0__pin_I01_1_, top_width_0_height_1_subtile_0__pin_I01_2_, top_width_0_height_1_subtile_0__pin_I01_3_, top_width_0_height_1_subtile_0__pin_I01_4_, top_width_0_height_1_subtile_0__pin_I01_5_, top_width_0_height_1_subtile_0__pin_I01_6_, top_width_0_height_1_subtile_0__pin_I01_7_, top_width_0_height_1_subtile_0__pin_I01_8_, top_width_0_height_1_subtile_0__pin_I01_9_, top_width_0_height_1_subtile_0__pin_I01_10_, top_width_0_height_1_subtile_0__pin_I01_11_}),
		.dsp_I11({top_width_0_height_1_subtile_0__pin_I11_0_, top_width_0_height_1_subtile_0__pin_I11_1_, top_width_0_height_1_subtile_0__pin_I11_2_, top_width_0_height_1_subtile_0__pin_I11_3_, top_width_0_height_1_subtile_0__pin_I11_4_, top_width_0_height_1_subtile_0__pin_I11_5_, top_width_0_height_1_subtile_0__pin_I11_6_, top_width_0_height_1_subtile_0__pin_I11_7_, top_width_0_height_1_subtile_0__pin_I11_8_, top_width_0_height_1_subtile_0__pin_I11_9_, top_width_0_height_1_subtile_0__pin_I11_10_, top_width_0_height_1_subtile_0__pin_I11_11_}),
		.dsp_I21({right_width_0_height_1_subtile_0__pin_I21_0_, right_width_0_height_1_subtile_0__pin_I21_1_, right_width_0_height_1_subtile_0__pin_I21_2_, right_width_0_height_1_subtile_0__pin_I21_3_, right_width_0_height_1_subtile_0__pin_I21_4_, right_width_0_height_1_subtile_0__pin_I21_5_, right_width_0_height_1_subtile_0__pin_I21_6_, right_width_0_height_1_subtile_0__pin_I21_7_, right_width_0_height_1_subtile_0__pin_I21_8_, right_width_0_height_1_subtile_0__pin_I21_9_, right_width_0_height_1_subtile_0__pin_I21_10_, right_width_0_height_1_subtile_0__pin_I21_11_}),
		.dsp_I31({right_width_0_height_1_subtile_0__pin_I31_0_, right_width_0_height_1_subtile_0__pin_I31_1_, right_width_0_height_1_subtile_0__pin_I31_2_, right_width_0_height_1_subtile_0__pin_I31_3_, right_width_0_height_1_subtile_0__pin_I31_4_, right_width_0_height_1_subtile_0__pin_I31_5_, right_width_0_height_1_subtile_0__pin_I31_6_, right_width_0_height_1_subtile_0__pin_I31_7_, right_width_0_height_1_subtile_0__pin_I31_8_, right_width_0_height_1_subtile_0__pin_I31_9_, right_width_0_height_1_subtile_0__pin_I31_10_, right_width_0_height_1_subtile_0__pin_I31_11_}),
		.dsp_IS1({top_width_0_height_1_subtile_0__pin_IS1_0_, top_width_0_height_1_subtile_0__pin_IS1_1_, top_width_0_height_1_subtile_0__pin_IS1_2_, right_width_0_height_1_subtile_0__pin_IS1_3_, right_width_0_height_1_subtile_0__pin_IS1_4_, right_width_0_height_1_subtile_0__pin_IS1_5_}),
		.dsp_I02({top_width_0_height_2_subtile_0__pin_I02_0_, top_width_0_height_2_subtile_0__pin_I02_1_, top_width_0_height_2_subtile_0__pin_I02_2_, top_width_0_height_2_subtile_0__pin_I02_3_, top_width_0_height_2_subtile_0__pin_I02_4_, top_width_0_height_2_subtile_0__pin_I02_5_, top_width_0_height_2_subtile_0__pin_I02_6_, top_width_0_height_2_subtile_0__pin_I02_7_, top_width_0_height_2_subtile_0__pin_I02_8_, top_width_0_height_2_subtile_0__pin_I02_9_, top_width_0_height_2_subtile_0__pin_I02_10_, top_width_0_height_2_subtile_0__pin_I02_11_}),
		.dsp_I12({top_width_0_height_2_subtile_0__pin_I12_0_, top_width_0_height_2_subtile_0__pin_I12_1_, top_width_0_height_2_subtile_0__pin_I12_2_, top_width_0_height_2_subtile_0__pin_I12_3_, top_width_0_height_2_subtile_0__pin_I12_4_, top_width_0_height_2_subtile_0__pin_I12_5_, top_width_0_height_2_subtile_0__pin_I12_6_, top_width_0_height_2_subtile_0__pin_I12_7_, top_width_0_height_2_subtile_0__pin_I12_8_, top_width_0_height_2_subtile_0__pin_I12_9_, top_width_0_height_2_subtile_0__pin_I12_10_, top_width_0_height_2_subtile_0__pin_I12_11_}),
		.dsp_I22({right_width_0_height_2_subtile_0__pin_I22_0_, right_width_0_height_2_subtile_0__pin_I22_1_, right_width_0_height_2_subtile_0__pin_I22_2_, right_width_0_height_2_subtile_0__pin_I22_3_, right_width_0_height_2_subtile_0__pin_I22_4_, right_width_0_height_2_subtile_0__pin_I22_5_, right_width_0_height_2_subtile_0__pin_I22_6_, right_width_0_height_2_subtile_0__pin_I22_7_, right_width_0_height_2_subtile_0__pin_I22_8_, right_width_0_height_2_subtile_0__pin_I22_9_, right_width_0_height_2_subtile_0__pin_I22_10_, right_width_0_height_2_subtile_0__pin_I22_11_}),
		.dsp_I32({right_width_0_height_2_subtile_0__pin_I32_0_, right_width_0_height_2_subtile_0__pin_I32_1_, right_width_0_height_2_subtile_0__pin_I32_2_, right_width_0_height_2_subtile_0__pin_I32_3_, right_width_0_height_2_subtile_0__pin_I32_4_, right_width_0_height_2_subtile_0__pin_I32_5_, right_width_0_height_2_subtile_0__pin_I32_6_, right_width_0_height_2_subtile_0__pin_I32_7_, right_width_0_height_2_subtile_0__pin_I32_8_, right_width_0_height_2_subtile_0__pin_I32_9_, right_width_0_height_2_subtile_0__pin_I32_10_, right_width_0_height_2_subtile_0__pin_I32_11_}),
		.dsp_IS2({top_width_0_height_2_subtile_0__pin_IS2_0_, top_width_0_height_2_subtile_0__pin_IS2_1_, top_width_0_height_2_subtile_0__pin_IS2_2_, right_width_0_height_2_subtile_0__pin_IS2_3_, right_width_0_height_2_subtile_0__pin_IS2_4_, right_width_0_height_2_subtile_0__pin_IS2_5_}),
		.dsp_sc_in({left_width_0_height_0_subtile_0__pin_sc_in_0_, left_width_0_height_0_subtile_0__pin_sc_in_1_, left_width_0_height_0_subtile_0__pin_sc_in_2_, left_width_0_height_0_subtile_0__pin_sc_in_3_, left_width_0_height_0_subtile_0__pin_sc_in_4_, left_width_0_height_0_subtile_0__pin_sc_in_5_, left_width_0_height_0_subtile_0__pin_sc_in_6_, left_width_0_height_0_subtile_0__pin_sc_in_7_, left_width_0_height_0_subtile_0__pin_sc_in_8_, left_width_0_height_0_subtile_0__pin_sc_in_9_, left_width_0_height_0_subtile_0__pin_sc_in_10_, left_width_0_height_0_subtile_0__pin_sc_in_11_, left_width_0_height_0_subtile_0__pin_sc_in_12_, left_width_0_height_0_subtile_0__pin_sc_in_13_, left_width_0_height_0_subtile_0__pin_sc_in_14_, left_width_0_height_0_subtile_0__pin_sc_in_15_, left_width_0_height_0_subtile_0__pin_sc_in_16_, left_width_0_height_0_subtile_0__pin_sc_in_17_, left_width_0_height_0_subtile_0__pin_sc_in_18_, left_width_0_height_0_subtile_0__pin_sc_in_19_}),
		.dsp_clk({left_width_0_height_0_subtile_0__pin_clk_0_, left_width_0_height_0_subtile_0__pin_clk_1_, left_width_0_height_0_subtile_0__pin_clk_2_, left_width_0_height_0_subtile_0__pin_clk_3_, left_width_0_height_0_subtile_0__pin_clk_4_, left_width_0_height_0_subtile_0__pin_clk_5_, left_width_0_height_0_subtile_0__pin_clk_6_, left_width_0_height_0_subtile_0__pin_clk_7_, left_width_0_height_0_subtile_0__pin_clk_8_, left_width_0_height_0_subtile_0__pin_clk_9_, left_width_0_height_0_subtile_0__pin_clk_10_, left_width_0_height_0_subtile_0__pin_clk_11_, left_width_0_height_0_subtile_0__pin_clk_12_, left_width_0_height_0_subtile_0__pin_clk_13_, left_width_0_height_0_subtile_0__pin_clk_14_, left_width_0_height_0_subtile_0__pin_clk_15_}),
		.ccff_head(ccff_head),
		.dsp_O0({top_width_0_height_0_subtile_0__pin_O0_0_, top_width_0_height_0_subtile_0__pin_O0_1_, top_width_0_height_0_subtile_0__pin_O0_2_, top_width_0_height_0_subtile_0__pin_O0_3_, top_width_0_height_0_subtile_0__pin_O0_4_, top_width_0_height_0_subtile_0__pin_O0_5_, top_width_0_height_0_subtile_0__pin_O0_6_, top_width_0_height_0_subtile_0__pin_O0_7_, top_width_0_height_0_subtile_0__pin_O0_8_, top_width_0_height_0_subtile_0__pin_O0_9_, top_width_0_height_0_subtile_0__pin_O0_10_, top_width_0_height_0_subtile_0__pin_O0_11_, right_width_0_height_0_subtile_0__pin_O0_12_, right_width_0_height_0_subtile_0__pin_O0_13_, right_width_0_height_0_subtile_0__pin_O0_14_, right_width_0_height_0_subtile_0__pin_O0_15_, right_width_0_height_0_subtile_0__pin_O0_16_, right_width_0_height_0_subtile_0__pin_O0_17_, right_width_0_height_0_subtile_0__pin_O0_18_, right_width_0_height_0_subtile_0__pin_O0_19_, right_width_0_height_0_subtile_0__pin_O0_20_, right_width_0_height_0_subtile_0__pin_O0_21_, right_width_0_height_0_subtile_0__pin_O0_22_, right_width_0_height_0_subtile_0__pin_O0_23_}),
		.dsp_O1({top_width_0_height_1_subtile_0__pin_O1_0_, top_width_0_height_1_subtile_0__pin_O1_1_, top_width_0_height_1_subtile_0__pin_O1_2_, top_width_0_height_1_subtile_0__pin_O1_3_, top_width_0_height_1_subtile_0__pin_O1_4_, top_width_0_height_1_subtile_0__pin_O1_5_, top_width_0_height_1_subtile_0__pin_O1_6_, top_width_0_height_1_subtile_0__pin_O1_7_, top_width_0_height_1_subtile_0__pin_O1_8_, top_width_0_height_1_subtile_0__pin_O1_9_, top_width_0_height_1_subtile_0__pin_O1_10_, top_width_0_height_1_subtile_0__pin_O1_11_, right_width_0_height_1_subtile_0__pin_O1_12_, right_width_0_height_1_subtile_0__pin_O1_13_, right_width_0_height_1_subtile_0__pin_O1_14_, right_width_0_height_1_subtile_0__pin_O1_15_, right_width_0_height_1_subtile_0__pin_O1_16_, right_width_0_height_1_subtile_0__pin_O1_17_, right_width_0_height_1_subtile_0__pin_O1_18_, right_width_0_height_1_subtile_0__pin_O1_19_, right_width_0_height_1_subtile_0__pin_O1_20_, right_width_0_height_1_subtile_0__pin_O1_21_, right_width_0_height_1_subtile_0__pin_O1_22_, right_width_0_height_1_subtile_0__pin_O1_23_}),
		.dsp_O2({top_width_0_height_2_subtile_0__pin_O2_0_, top_width_0_height_2_subtile_0__pin_O2_1_, top_width_0_height_2_subtile_0__pin_O2_2_, top_width_0_height_2_subtile_0__pin_O2_3_, top_width_0_height_2_subtile_0__pin_O2_4_, top_width_0_height_2_subtile_0__pin_O2_5_, top_width_0_height_2_subtile_0__pin_O2_6_, top_width_0_height_2_subtile_0__pin_O2_7_, top_width_0_height_2_subtile_0__pin_O2_8_, top_width_0_height_2_subtile_0__pin_O2_9_, top_width_0_height_2_subtile_0__pin_O2_10_, top_width_0_height_2_subtile_0__pin_O2_11_, right_width_0_height_2_subtile_0__pin_O2_12_, right_width_0_height_2_subtile_0__pin_O2_13_, right_width_0_height_2_subtile_0__pin_O2_14_, right_width_0_height_2_subtile_0__pin_O2_15_, right_width_0_height_2_subtile_0__pin_O2_16_, right_width_0_height_2_subtile_0__pin_O2_17_, right_width_0_height_2_subtile_0__pin_O2_18_, right_width_0_height_2_subtile_0__pin_O2_19_, right_width_0_height_2_subtile_0__pin_O2_20_, right_width_0_height_2_subtile_0__pin_O2_21_, right_width_0_height_2_subtile_0__pin_O2_22_, right_width_0_height_2_subtile_0__pin_O2_23_}),
		.dsp_sc_out({right_width_0_height_0_subtile_0__pin_sc_out_0_, right_width_0_height_0_subtile_0__pin_sc_out_1_, right_width_0_height_0_subtile_0__pin_sc_out_2_, right_width_0_height_0_subtile_0__pin_sc_out_3_, right_width_0_height_0_subtile_0__pin_sc_out_4_, right_width_0_height_0_subtile_0__pin_sc_out_5_, right_width_0_height_0_subtile_0__pin_sc_out_6_, right_width_0_height_0_subtile_0__pin_sc_out_7_, right_width_0_height_0_subtile_0__pin_sc_out_8_, right_width_0_height_0_subtile_0__pin_sc_out_9_, right_width_0_height_0_subtile_0__pin_sc_out_10_, right_width_0_height_0_subtile_0__pin_sc_out_11_, right_width_0_height_0_subtile_0__pin_sc_out_12_, right_width_0_height_0_subtile_0__pin_sc_out_13_, right_width_0_height_0_subtile_0__pin_sc_out_14_, right_width_0_height_0_subtile_0__pin_sc_out_15_, right_width_0_height_0_subtile_0__pin_sc_out_16_, right_width_0_height_0_subtile_0__pin_sc_out_17_, right_width_0_height_0_subtile_0__pin_sc_out_18_, right_width_0_height_0_subtile_0__pin_sc_out_19_}),
		.ccff_tail(ccff_tail));

endmodule
// ----- END Verilog module for grid_dsp -----

//----- Default net type -----
`default_nettype none



// ----- END Grid Verilog module: grid_dsp -----

