//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for Unique Switch Blocks[2][8]
//	Author: Xifan TANG
//	Organization: University of Utah
//-------------------------------------------
//----- Time scale -----
`timescale 1ns / 1ps

//----- Default net type -----
`default_nettype wire

// ----- Verilog module for sb_2__8_ -----
module sb_2__8_(config_enable,
                prog_clock,
                chanx_right_in,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_8__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_9__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_10__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_11__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_24__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_25__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_26__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_27__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_28__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_29__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_30__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_31__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_32__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_33__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_34__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_35__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_36__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_37__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_38__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_39__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_40__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_41__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_42__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_43__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_44__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_45__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_46__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_47__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_48__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_49__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_50__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_51__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_52__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_53__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_54__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_55__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_56__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_57__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_58__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_59__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_60__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_61__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_62__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_63__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_64__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_65__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_66__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_67__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_68__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_69__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_70__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_71__pin_a2f_o_0_,
                chany_bottom_in,
                bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_,
                bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_,
                bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_,
                bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_,
                bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_,
                bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_,
                bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_,
                bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_,
                bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_,
                bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_,
                bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_,
                bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_,
                chanx_left_in,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_8__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_9__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_10__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_11__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_24__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_25__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_26__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_27__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_28__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_29__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_30__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_31__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_32__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_33__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_34__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_35__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_36__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_37__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_38__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_39__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_40__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_41__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_42__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_43__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_44__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_45__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_46__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_47__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_48__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_49__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_50__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_51__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_52__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_53__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_54__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_55__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_56__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_57__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_58__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_59__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_60__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_61__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_62__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_63__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_64__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_65__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_66__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_67__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_68__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_69__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_70__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_71__pin_a2f_o_0_,
                ccff_head,
                chanx_right_out,
                chany_bottom_out,
                chanx_left_out,
                ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_clock;
//----- INPUT PORTS -----
input [0:95] chanx_right_in;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_8__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_9__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_10__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_11__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_24__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_25__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_26__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_27__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_28__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_29__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_30__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_31__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_32__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_33__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_34__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_35__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_36__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_37__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_38__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_39__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_40__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_41__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_42__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_43__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_44__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_45__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_46__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_47__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_48__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_49__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_50__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_51__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_52__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_53__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_54__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_55__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_56__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_57__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_58__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_59__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_60__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_61__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_62__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_63__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_64__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_65__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_66__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_67__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_68__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_69__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_70__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_71__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:95] chany_bottom_in;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:95] chanx_left_in;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_8__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_9__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_10__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_11__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_24__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_25__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_26__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_27__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_28__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_29__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_30__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_31__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_32__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_33__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_34__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_35__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_36__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_37__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_38__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_39__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_40__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_41__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_42__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_43__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_44__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_45__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_46__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_47__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_48__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_49__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_50__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_51__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_52__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_53__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_54__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_55__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_56__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_57__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_58__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_59__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_60__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_61__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_62__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_63__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_64__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_65__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_66__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_67__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_68__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_69__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_70__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_71__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:95] chanx_right_out;
//----- OUTPUT PORTS -----
output [0:95] chany_bottom_out;
//----- OUTPUT PORTS -----
output [0:95] chanx_left_out;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:3] mux_tree_tapbuf_L2SB_size11_0_sram;
wire [0:3] mux_tree_tapbuf_L2SB_size11_0_sram_inv;
wire [0:3] mux_tree_tapbuf_L2SB_size11_1_sram;
wire [0:3] mux_tree_tapbuf_L2SB_size11_1_sram_inv;
wire [0:3] mux_tree_tapbuf_L2SB_size11_2_sram;
wire [0:3] mux_tree_tapbuf_L2SB_size11_2_sram_inv;
wire [0:3] mux_tree_tapbuf_L2SB_size11_3_sram;
wire [0:3] mux_tree_tapbuf_L2SB_size11_3_sram_inv;
wire [0:3] mux_tree_tapbuf_L2SB_size11_4_sram;
wire [0:3] mux_tree_tapbuf_L2SB_size11_4_sram_inv;
wire [0:3] mux_tree_tapbuf_L2SB_size11_5_sram;
wire [0:3] mux_tree_tapbuf_L2SB_size11_5_sram_inv;
wire [0:3] mux_tree_tapbuf_L2SB_size11_6_sram;
wire [0:3] mux_tree_tapbuf_L2SB_size11_6_sram_inv;
wire [0:3] mux_tree_tapbuf_L2SB_size12_0_sram;
wire [0:3] mux_tree_tapbuf_L2SB_size12_0_sram_inv;
wire [0:3] mux_tree_tapbuf_L2SB_size12_1_sram;
wire [0:3] mux_tree_tapbuf_L2SB_size12_1_sram_inv;
wire [0:3] mux_tree_tapbuf_L2SB_size12_2_sram;
wire [0:3] mux_tree_tapbuf_L2SB_size12_2_sram_inv;
wire [0:3] mux_tree_tapbuf_L2SB_size12_3_sram;
wire [0:3] mux_tree_tapbuf_L2SB_size12_3_sram_inv;
wire [0:3] mux_tree_tapbuf_L2SB_size12_4_sram;
wire [0:3] mux_tree_tapbuf_L2SB_size12_4_sram_inv;
wire [0:3] mux_tree_tapbuf_L2SB_size12_5_sram;
wire [0:3] mux_tree_tapbuf_L2SB_size12_5_sram_inv;
wire [0:3] mux_tree_tapbuf_L2SB_size12_6_sram;
wire [0:3] mux_tree_tapbuf_L2SB_size12_6_sram_inv;
wire [0:3] mux_tree_tapbuf_L2SB_size12_7_sram;
wire [0:3] mux_tree_tapbuf_L2SB_size12_7_sram_inv;
wire [0:3] mux_tree_tapbuf_L2SB_size13_0_sram;
wire [0:3] mux_tree_tapbuf_L2SB_size13_0_sram_inv;
wire [0:3] mux_tree_tapbuf_L2SB_size13_1_sram;
wire [0:3] mux_tree_tapbuf_L2SB_size13_1_sram_inv;
wire [0:3] mux_tree_tapbuf_L2SB_size13_2_sram;
wire [0:3] mux_tree_tapbuf_L2SB_size13_2_sram_inv;
wire [0:3] mux_tree_tapbuf_L2SB_size13_3_sram;
wire [0:3] mux_tree_tapbuf_L2SB_size13_3_sram_inv;
wire [0:3] mux_tree_tapbuf_L2SB_size13_4_sram;
wire [0:3] mux_tree_tapbuf_L2SB_size13_4_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size3_0_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size3_0_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size3_1_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size3_1_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size3_2_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size3_2_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size3_3_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size3_3_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size3_4_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size3_4_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size3_5_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size3_5_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size3_6_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size3_6_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_0_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_0_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_10_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_10_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_11_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_11_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_1_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_1_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_2_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_2_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_3_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_3_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_4_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_4_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_5_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_5_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_6_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_6_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_7_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_7_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_8_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_8_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_9_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_9_sram_inv;
wire [0:4] mux_tree_tapbuf_L4SB_size17_0_sram;
wire [0:4] mux_tree_tapbuf_L4SB_size17_0_sram_inv;
wire [0:4] mux_tree_tapbuf_L4SB_size17_10_sram;
wire [0:4] mux_tree_tapbuf_L4SB_size17_10_sram_inv;
wire [0:4] mux_tree_tapbuf_L4SB_size17_11_sram;
wire [0:4] mux_tree_tapbuf_L4SB_size17_11_sram_inv;
wire [0:4] mux_tree_tapbuf_L4SB_size17_12_sram;
wire [0:4] mux_tree_tapbuf_L4SB_size17_12_sram_inv;
wire [0:4] mux_tree_tapbuf_L4SB_size17_13_sram;
wire [0:4] mux_tree_tapbuf_L4SB_size17_13_sram_inv;
wire [0:4] mux_tree_tapbuf_L4SB_size17_14_sram;
wire [0:4] mux_tree_tapbuf_L4SB_size17_14_sram_inv;
wire [0:4] mux_tree_tapbuf_L4SB_size17_15_sram;
wire [0:4] mux_tree_tapbuf_L4SB_size17_15_sram_inv;
wire [0:4] mux_tree_tapbuf_L4SB_size17_16_sram;
wire [0:4] mux_tree_tapbuf_L4SB_size17_16_sram_inv;
wire [0:4] mux_tree_tapbuf_L4SB_size17_17_sram;
wire [0:4] mux_tree_tapbuf_L4SB_size17_17_sram_inv;
wire [0:4] mux_tree_tapbuf_L4SB_size17_18_sram;
wire [0:4] mux_tree_tapbuf_L4SB_size17_18_sram_inv;
wire [0:4] mux_tree_tapbuf_L4SB_size17_19_sram;
wire [0:4] mux_tree_tapbuf_L4SB_size17_19_sram_inv;
wire [0:4] mux_tree_tapbuf_L4SB_size17_1_sram;
wire [0:4] mux_tree_tapbuf_L4SB_size17_1_sram_inv;
wire [0:4] mux_tree_tapbuf_L4SB_size17_20_sram;
wire [0:4] mux_tree_tapbuf_L4SB_size17_20_sram_inv;
wire [0:4] mux_tree_tapbuf_L4SB_size17_21_sram;
wire [0:4] mux_tree_tapbuf_L4SB_size17_21_sram_inv;
wire [0:4] mux_tree_tapbuf_L4SB_size17_22_sram;
wire [0:4] mux_tree_tapbuf_L4SB_size17_22_sram_inv;
wire [0:4] mux_tree_tapbuf_L4SB_size17_23_sram;
wire [0:4] mux_tree_tapbuf_L4SB_size17_23_sram_inv;
wire [0:4] mux_tree_tapbuf_L4SB_size17_24_sram;
wire [0:4] mux_tree_tapbuf_L4SB_size17_24_sram_inv;
wire [0:4] mux_tree_tapbuf_L4SB_size17_25_sram;
wire [0:4] mux_tree_tapbuf_L4SB_size17_25_sram_inv;
wire [0:4] mux_tree_tapbuf_L4SB_size17_26_sram;
wire [0:4] mux_tree_tapbuf_L4SB_size17_26_sram_inv;
wire [0:4] mux_tree_tapbuf_L4SB_size17_27_sram;
wire [0:4] mux_tree_tapbuf_L4SB_size17_27_sram_inv;
wire [0:4] mux_tree_tapbuf_L4SB_size17_28_sram;
wire [0:4] mux_tree_tapbuf_L4SB_size17_28_sram_inv;
wire [0:4] mux_tree_tapbuf_L4SB_size17_29_sram;
wire [0:4] mux_tree_tapbuf_L4SB_size17_29_sram_inv;
wire [0:4] mux_tree_tapbuf_L4SB_size17_2_sram;
wire [0:4] mux_tree_tapbuf_L4SB_size17_2_sram_inv;
wire [0:4] mux_tree_tapbuf_L4SB_size17_30_sram;
wire [0:4] mux_tree_tapbuf_L4SB_size17_30_sram_inv;
wire [0:4] mux_tree_tapbuf_L4SB_size17_31_sram;
wire [0:4] mux_tree_tapbuf_L4SB_size17_31_sram_inv;
wire [0:4] mux_tree_tapbuf_L4SB_size17_32_sram;
wire [0:4] mux_tree_tapbuf_L4SB_size17_32_sram_inv;
wire [0:4] mux_tree_tapbuf_L4SB_size17_33_sram;
wire [0:4] mux_tree_tapbuf_L4SB_size17_33_sram_inv;
wire [0:4] mux_tree_tapbuf_L4SB_size17_3_sram;
wire [0:4] mux_tree_tapbuf_L4SB_size17_3_sram_inv;
wire [0:4] mux_tree_tapbuf_L4SB_size17_4_sram;
wire [0:4] mux_tree_tapbuf_L4SB_size17_4_sram_inv;
wire [0:4] mux_tree_tapbuf_L4SB_size17_5_sram;
wire [0:4] mux_tree_tapbuf_L4SB_size17_5_sram_inv;
wire [0:4] mux_tree_tapbuf_L4SB_size17_6_sram;
wire [0:4] mux_tree_tapbuf_L4SB_size17_6_sram_inv;
wire [0:4] mux_tree_tapbuf_L4SB_size17_7_sram;
wire [0:4] mux_tree_tapbuf_L4SB_size17_7_sram_inv;
wire [0:4] mux_tree_tapbuf_L4SB_size17_8_sram;
wire [0:4] mux_tree_tapbuf_L4SB_size17_8_sram_inv;
wire [0:4] mux_tree_tapbuf_L4SB_size17_9_sram;
wire [0:4] mux_tree_tapbuf_L4SB_size17_9_sram_inv;
wire [0:4] mux_tree_tapbuf_L4SB_size18_0_sram;
wire [0:4] mux_tree_tapbuf_L4SB_size18_0_sram_inv;
wire [0:4] mux_tree_tapbuf_L4SB_size18_1_sram;
wire [0:4] mux_tree_tapbuf_L4SB_size18_1_sram_inv;
wire [0:4] mux_tree_tapbuf_L4SB_size18_2_sram;
wire [0:4] mux_tree_tapbuf_L4SB_size18_2_sram_inv;
wire [0:4] mux_tree_tapbuf_L4SB_size18_3_sram;
wire [0:4] mux_tree_tapbuf_L4SB_size18_3_sram_inv;
wire [0:4] mux_tree_tapbuf_L4SB_size18_4_sram;
wire [0:4] mux_tree_tapbuf_L4SB_size18_4_sram_inv;
wire [0:4] mux_tree_tapbuf_L4SB_size18_5_sram;
wire [0:4] mux_tree_tapbuf_L4SB_size18_5_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_0_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_0_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_10_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_10_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_11_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_11_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_12_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_12_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_13_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_13_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_14_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_14_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_15_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_15_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_16_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_16_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_17_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_17_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_18_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_18_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_19_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_19_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_1_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_1_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_20_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_20_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_21_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_21_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_22_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_22_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_23_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_23_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_24_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_24_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_25_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_25_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_26_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_26_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_27_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_27_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_28_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_28_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_29_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_29_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_2_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_2_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_3_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_3_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_4_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_4_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_5_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_5_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_6_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_6_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_7_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_7_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_8_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_8_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_9_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_9_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_0_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_0_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_10_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_10_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_11_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_11_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_12_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_12_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_13_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_13_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_14_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_14_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_15_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_15_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_16_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_16_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_17_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_17_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_18_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_18_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_19_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_19_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_1_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_1_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_20_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_20_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_21_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_21_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_22_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_22_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_23_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_23_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_24_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_24_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_25_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_25_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_26_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_26_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_27_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_27_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_2_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_2_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_3_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_3_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_4_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_4_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_5_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_5_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_6_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_6_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_7_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_7_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_8_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_8_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_9_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_9_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_0_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_0_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_1_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_1_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_2_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_2_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_3_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_3_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_4_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_4_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_5_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_5_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_6_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_6_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_7_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_7_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_8_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_8_sram_inv;

// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[1] = chanx_right_in[0];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[3] = chanx_right_in[2];
// ----- Local connection due to Wire 4 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[5] = chanx_right_in[4];
// ----- Local connection due to Wire 6 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[7] = chanx_right_in[6];
// ----- Local connection due to Wire 8 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[9] = chanx_right_in[8];
// ----- Local connection due to Wire 10 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[11] = chanx_right_in[10];
// ----- Local connection due to Wire 12 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[13] = chanx_right_in[12];
// ----- Local connection due to Wire 14 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[15] = chanx_right_in[14];
// ----- Local connection due to Wire 16 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[17] = chanx_right_in[16];
// ----- Local connection due to Wire 19 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[20] = chanx_right_in[19];
// ----- Local connection due to Wire 20 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[21] = chanx_right_in[20];
// ----- Local connection due to Wire 21 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[22] = chanx_right_in[21];
// ----- Local connection due to Wire 23 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[24] = chanx_right_in[23];
// ----- Local connection due to Wire 24 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[25] = chanx_right_in[24];
// ----- Local connection due to Wire 25 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[26] = chanx_right_in[25];
// ----- Local connection due to Wire 27 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[28] = chanx_right_in[27];
// ----- Local connection due to Wire 28 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[29] = chanx_right_in[28];
// ----- Local connection due to Wire 29 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[30] = chanx_right_in[29];
// ----- Local connection due to Wire 31 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[32] = chanx_right_in[31];
// ----- Local connection due to Wire 32 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[33] = chanx_right_in[32];
// ----- Local connection due to Wire 33 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[34] = chanx_right_in[33];
// ----- Local connection due to Wire 35 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[36] = chanx_right_in[35];
// ----- Local connection due to Wire 36 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[37] = chanx_right_in[36];
// ----- Local connection due to Wire 37 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[38] = chanx_right_in[37];
// ----- Local connection due to Wire 39 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[40] = chanx_right_in[39];
// ----- Local connection due to Wire 40 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[41] = chanx_right_in[40];
// ----- Local connection due to Wire 41 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[42] = chanx_right_in[41];
// ----- Local connection due to Wire 43 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[44] = chanx_right_in[43];
// ----- Local connection due to Wire 44 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[45] = chanx_right_in[44];
// ----- Local connection due to Wire 45 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[46] = chanx_right_in[45];
// ----- Local connection due to Wire 47 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[48] = chanx_right_in[47];
// ----- Local connection due to Wire 48 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[49] = chanx_right_in[48];
// ----- Local connection due to Wire 49 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[50] = chanx_right_in[49];
// ----- Local connection due to Wire 51 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[52] = chanx_right_in[51];
// ----- Local connection due to Wire 52 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[53] = chanx_right_in[52];
// ----- Local connection due to Wire 53 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[54] = chanx_right_in[53];
// ----- Local connection due to Wire 55 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[56] = chanx_right_in[55];
// ----- Local connection due to Wire 56 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[57] = chanx_right_in[56];
// ----- Local connection due to Wire 57 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[58] = chanx_right_in[57];
// ----- Local connection due to Wire 59 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[60] = chanx_right_in[59];
// ----- Local connection due to Wire 60 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[61] = chanx_right_in[60];
// ----- Local connection due to Wire 61 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[62] = chanx_right_in[61];
// ----- Local connection due to Wire 63 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[64] = chanx_right_in[63];
// ----- Local connection due to Wire 64 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[65] = chanx_right_in[64];
// ----- Local connection due to Wire 65 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[66] = chanx_right_in[65];
// ----- Local connection due to Wire 67 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[68] = chanx_right_in[67];
// ----- Local connection due to Wire 68 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[69] = chanx_right_in[68];
// ----- Local connection due to Wire 69 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[70] = chanx_right_in[69];
// ----- Local connection due to Wire 71 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[72] = chanx_right_in[71];
// ----- Local connection due to Wire 72 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[73] = chanx_right_in[72];
// ----- Local connection due to Wire 73 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[74] = chanx_right_in[73];
// ----- Local connection due to Wire 75 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[76] = chanx_right_in[75];
// ----- Local connection due to Wire 76 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[77] = chanx_right_in[76];
// ----- Local connection due to Wire 77 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[78] = chanx_right_in[77];
// ----- Local connection due to Wire 79 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[80] = chanx_right_in[79];
// ----- Local connection due to Wire 80 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[81] = chanx_right_in[80];
// ----- Local connection due to Wire 81 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[82] = chanx_right_in[81];
// ----- Local connection due to Wire 83 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[84] = chanx_right_in[83];
// ----- Local connection due to Wire 84 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[85] = chanx_right_in[84];
// ----- Local connection due to Wire 85 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[86] = chanx_right_in[85];
// ----- Local connection due to Wire 87 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[88] = chanx_right_in[87];
// ----- Local connection due to Wire 88 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[89] = chanx_right_in[88];
// ----- Local connection due to Wire 89 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[90] = chanx_right_in[89];
// ----- Local connection due to Wire 91 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[92] = chanx_right_in[91];
// ----- Local connection due to Wire 92 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[93] = chanx_right_in[92];
// ----- Local connection due to Wire 93 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[94] = chanx_right_in[93];
// ----- Local connection due to Wire 264 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[1] = chanx_left_in[0];
// ----- Local connection due to Wire 266 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[3] = chanx_left_in[2];
// ----- Local connection due to Wire 268 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[5] = chanx_left_in[4];
// ----- Local connection due to Wire 270 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[7] = chanx_left_in[6];
// ----- Local connection due to Wire 272 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[9] = chanx_left_in[8];
// ----- Local connection due to Wire 274 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[11] = chanx_left_in[10];
// ----- Local connection due to Wire 276 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[13] = chanx_left_in[12];
// ----- Local connection due to Wire 278 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[15] = chanx_left_in[14];
// ----- Local connection due to Wire 280 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[17] = chanx_left_in[16];
// ----- Local connection due to Wire 283 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[20] = chanx_left_in[19];
// ----- Local connection due to Wire 284 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[21] = chanx_left_in[20];
// ----- Local connection due to Wire 285 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[22] = chanx_left_in[21];
// ----- Local connection due to Wire 287 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[24] = chanx_left_in[23];
// ----- Local connection due to Wire 288 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[25] = chanx_left_in[24];
// ----- Local connection due to Wire 289 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[26] = chanx_left_in[25];
// ----- Local connection due to Wire 291 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[28] = chanx_left_in[27];
// ----- Local connection due to Wire 292 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[29] = chanx_left_in[28];
// ----- Local connection due to Wire 293 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[30] = chanx_left_in[29];
// ----- Local connection due to Wire 295 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[32] = chanx_left_in[31];
// ----- Local connection due to Wire 296 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[33] = chanx_left_in[32];
// ----- Local connection due to Wire 297 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[34] = chanx_left_in[33];
// ----- Local connection due to Wire 299 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[36] = chanx_left_in[35];
// ----- Local connection due to Wire 300 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[37] = chanx_left_in[36];
// ----- Local connection due to Wire 301 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[38] = chanx_left_in[37];
// ----- Local connection due to Wire 303 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[40] = chanx_left_in[39];
// ----- Local connection due to Wire 304 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[41] = chanx_left_in[40];
// ----- Local connection due to Wire 305 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[42] = chanx_left_in[41];
// ----- Local connection due to Wire 307 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[44] = chanx_left_in[43];
// ----- Local connection due to Wire 308 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[45] = chanx_left_in[44];
// ----- Local connection due to Wire 309 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[46] = chanx_left_in[45];
// ----- Local connection due to Wire 311 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[48] = chanx_left_in[47];
// ----- Local connection due to Wire 312 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[49] = chanx_left_in[48];
// ----- Local connection due to Wire 313 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[50] = chanx_left_in[49];
// ----- Local connection due to Wire 315 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[52] = chanx_left_in[51];
// ----- Local connection due to Wire 316 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[53] = chanx_left_in[52];
// ----- Local connection due to Wire 317 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[54] = chanx_left_in[53];
// ----- Local connection due to Wire 319 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[56] = chanx_left_in[55];
// ----- Local connection due to Wire 320 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[57] = chanx_left_in[56];
// ----- Local connection due to Wire 321 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[58] = chanx_left_in[57];
// ----- Local connection due to Wire 323 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[60] = chanx_left_in[59];
// ----- Local connection due to Wire 324 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[61] = chanx_left_in[60];
// ----- Local connection due to Wire 325 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[62] = chanx_left_in[61];
// ----- Local connection due to Wire 327 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[64] = chanx_left_in[63];
// ----- Local connection due to Wire 328 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[65] = chanx_left_in[64];
// ----- Local connection due to Wire 329 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[66] = chanx_left_in[65];
// ----- Local connection due to Wire 331 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[68] = chanx_left_in[67];
// ----- Local connection due to Wire 332 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[69] = chanx_left_in[68];
// ----- Local connection due to Wire 333 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[70] = chanx_left_in[69];
// ----- Local connection due to Wire 335 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[72] = chanx_left_in[71];
// ----- Local connection due to Wire 336 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[73] = chanx_left_in[72];
// ----- Local connection due to Wire 337 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[74] = chanx_left_in[73];
// ----- Local connection due to Wire 339 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[76] = chanx_left_in[75];
// ----- Local connection due to Wire 340 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[77] = chanx_left_in[76];
// ----- Local connection due to Wire 341 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[78] = chanx_left_in[77];
// ----- Local connection due to Wire 343 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[80] = chanx_left_in[79];
// ----- Local connection due to Wire 344 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[81] = chanx_left_in[80];
// ----- Local connection due to Wire 345 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[82] = chanx_left_in[81];
// ----- Local connection due to Wire 347 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[84] = chanx_left_in[83];
// ----- Local connection due to Wire 348 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[85] = chanx_left_in[84];
// ----- Local connection due to Wire 349 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[86] = chanx_left_in[85];
// ----- Local connection due to Wire 351 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[88] = chanx_left_in[87];
// ----- Local connection due to Wire 352 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[89] = chanx_left_in[88];
// ----- Local connection due to Wire 353 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[90] = chanx_left_in[89];
// ----- Local connection due to Wire 355 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[92] = chanx_left_in[91];
// ----- Local connection due to Wire 356 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[93] = chanx_left_in[92];
// ----- Local connection due to Wire 357 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[94] = chanx_left_in[93];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	mux_tree_tapbuf_L2SB_size12 mux_right_track_0 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_10__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_32__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_42__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_52__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_62__pin_a2f_o_0_, chany_bottom_in[28], chany_bottom_in[58], chany_bottom_in[88], chanx_left_in[0], chanx_left_in[47], chanx_left_in[87]}),
		.sram(mux_tree_tapbuf_L2SB_size12_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L2SB_size12_0_sram_inv[0:3]),
		.out(chanx_right_out[0]));

	mux_tree_tapbuf_L2SB_size12 mux_right_track_4 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_11__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_33__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_43__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_53__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_63__pin_a2f_o_0_, chany_bottom_in[27], chany_bottom_in[57], chany_bottom_in[87], chanx_left_in[2], chanx_left_in[48], chanx_left_in[88]}),
		.sram(mux_tree_tapbuf_L2SB_size12_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L2SB_size12_1_sram_inv[0:3]),
		.out(chanx_right_out[2]));

	mux_tree_tapbuf_L2SB_size12 mux_right_track_8 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_24__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_34__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_44__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_54__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_64__pin_a2f_o_0_, chany_bottom_in[26], chany_bottom_in[56], chany_bottom_in[86], chanx_left_in[4], chanx_left_in[49], chanx_left_in[89]}),
		.sram(mux_tree_tapbuf_L2SB_size12_2_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L2SB_size12_2_sram_inv[0:3]),
		.out(chanx_right_out[4]));

	mux_tree_tapbuf_L2SB_size12 mux_right_track_12 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_25__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_35__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_45__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_55__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_65__pin_a2f_o_0_, chany_bottom_in[25], chany_bottom_in[55], chany_bottom_in[85], chanx_left_in[6], chanx_left_in[51], chanx_left_in[91]}),
		.sram(mux_tree_tapbuf_L2SB_size12_3_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L2SB_size12_3_sram_inv[0:3]),
		.out(chanx_right_out[6]));

	mux_tree_tapbuf_L2SB_size12 mux_right_track_16 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_26__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_36__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_46__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_56__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_66__pin_a2f_o_0_, chany_bottom_in[24], chany_bottom_in[54], chany_bottom_in[84], chanx_left_in[8], chanx_left_in[52], chanx_left_in[92]}),
		.sram(mux_tree_tapbuf_L2SB_size12_4_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L2SB_size12_4_sram_inv[0:3]),
		.out(chanx_right_out[8]));

	mux_tree_tapbuf_L2SB_size12 mux_right_track_20 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_27__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_37__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_47__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_57__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_67__pin_a2f_o_0_, chany_bottom_in[23], chany_bottom_in[53], chany_bottom_in[83], chanx_left_in[10], chanx_left_in[53], chanx_left_in[93]}),
		.sram(mux_tree_tapbuf_L2SB_size12_5_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L2SB_size12_5_sram_inv[0:3]),
		.out(chanx_right_out[10]));

	mux_tree_tapbuf_L2SB_size12 mux_left_track_1 (
		.in({chanx_right_in[0], chanx_right_in[47], chanx_right_in[87], chany_bottom_in[29], chany_bottom_in[59], chany_bottom_in[89], left_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_10__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_32__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_42__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_52__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_62__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L2SB_size12_6_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L2SB_size12_6_sram_inv[0:3]),
		.out(chanx_left_out[0]));

	mux_tree_tapbuf_L2SB_size12 mux_left_track_25 (
		.in({chanx_right_in[12], chanx_right_in[55], chany_bottom_in[5], chany_bottom_in[35], chany_bottom_in[65], chany_bottom_in[95], left_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_28__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_38__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_48__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_58__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_68__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L2SB_size12_7_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L2SB_size12_7_sram_inv[0:3]),
		.out(chanx_left_out[12]));

	mux_tree_tapbuf_L2SB_size12_mem mem_right_track_0 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(ccff_head),
		.ccff_tail(mux_tree_tapbuf_L2SB_size12_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size12_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L2SB_size12_0_sram_inv[0:3]));

	mux_tree_tapbuf_L2SB_size12_mem mem_right_track_4 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size12_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size12_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size12_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L2SB_size12_1_sram_inv[0:3]));

	mux_tree_tapbuf_L2SB_size12_mem mem_right_track_8 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size12_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size12_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size12_2_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L2SB_size12_2_sram_inv[0:3]));

	mux_tree_tapbuf_L2SB_size12_mem mem_right_track_12 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size12_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size12_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size12_3_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L2SB_size12_3_sram_inv[0:3]));

	mux_tree_tapbuf_L2SB_size12_mem mem_right_track_16 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size12_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size12_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size12_4_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L2SB_size12_4_sram_inv[0:3]));

	mux_tree_tapbuf_L2SB_size12_mem mem_right_track_20 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size12_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size12_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size12_5_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L2SB_size12_5_sram_inv[0:3]));

	mux_tree_tapbuf_L2SB_size12_mem mem_left_track_1 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size2_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size12_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size12_6_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L2SB_size12_6_sram_inv[0:3]));

	mux_tree_tapbuf_L2SB_size12_mem mem_left_track_25 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size13_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size12_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size12_7_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L2SB_size12_7_sram_inv[0:3]));

	mux_tree_tapbuf_L2SB_size11 mux_right_track_24 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_28__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_38__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_48__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_58__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_68__pin_a2f_o_0_, chany_bottom_in[22], chany_bottom_in[52], chany_bottom_in[82], chanx_left_in[12], chanx_left_in[55]}),
		.sram(mux_tree_tapbuf_L2SB_size11_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L2SB_size11_0_sram_inv[0:3]),
		.out(chanx_right_out[12]));

	mux_tree_tapbuf_L2SB_size11 mux_right_track_28 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_29__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_39__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_49__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_59__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_69__pin_a2f_o_0_, chany_bottom_in[21], chany_bottom_in[51], chany_bottom_in[81], chanx_left_in[14], chanx_left_in[56]}),
		.sram(mux_tree_tapbuf_L2SB_size11_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L2SB_size11_1_sram_inv[0:3]),
		.out(chanx_right_out[14]));

	mux_tree_tapbuf_L2SB_size11 mux_right_track_32 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_8__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_30__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_40__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_50__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_60__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_70__pin_a2f_o_0_, chany_bottom_in[20], chany_bottom_in[50], chany_bottom_in[80], chanx_left_in[16], chanx_left_in[57]}),
		.sram(mux_tree_tapbuf_L2SB_size11_2_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L2SB_size11_2_sram_inv[0:3]),
		.out(chanx_right_out[16]));

	mux_tree_tapbuf_L2SB_size11 mux_right_track_36 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_9__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_31__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_41__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_51__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_61__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_71__pin_a2f_o_0_, chany_bottom_in[19], chany_bottom_in[49], chany_bottom_in[79], chanx_left_in[19], chanx_left_in[59]}),
		.sram(mux_tree_tapbuf_L2SB_size11_3_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L2SB_size11_3_sram_inv[0:3]),
		.out(chanx_right_out[18]));

	mux_tree_tapbuf_L2SB_size11 mux_left_track_29 (
		.in({chanx_right_in[14], chanx_right_in[56], chany_bottom_in[6], chany_bottom_in[36], chany_bottom_in[66], left_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_29__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_39__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_49__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_59__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_69__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L2SB_size11_4_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L2SB_size11_4_sram_inv[0:3]),
		.out(chanx_left_out[14]));

	mux_tree_tapbuf_L2SB_size11 mux_left_track_33 (
		.in({chanx_right_in[16], chanx_right_in[57], chany_bottom_in[7], chany_bottom_in[37], chany_bottom_in[67], left_bottom_grid_top_width_0_height_0_subtile_8__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_30__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_40__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_50__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_60__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_70__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L2SB_size11_5_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L2SB_size11_5_sram_inv[0:3]),
		.out(chanx_left_out[16]));

	mux_tree_tapbuf_L2SB_size11 mux_left_track_37 (
		.in({chanx_right_in[19], chanx_right_in[59], chany_bottom_in[8], chany_bottom_in[38], chany_bottom_in[68], left_bottom_grid_top_width_0_height_0_subtile_9__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_31__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_41__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_51__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_61__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_71__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L2SB_size11_6_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L2SB_size11_6_sram_inv[0:3]),
		.out(chanx_left_out[18]));

	mux_tree_tapbuf_L2SB_size11_mem mem_right_track_24 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size12_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size11_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size11_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L2SB_size11_0_sram_inv[0:3]));

	mux_tree_tapbuf_L2SB_size11_mem mem_right_track_28 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size11_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size11_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size11_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L2SB_size11_1_sram_inv[0:3]));

	mux_tree_tapbuf_L2SB_size11_mem mem_right_track_32 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size11_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size11_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size11_2_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L2SB_size11_2_sram_inv[0:3]));

	mux_tree_tapbuf_L2SB_size11_mem mem_right_track_36 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size11_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size11_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size11_3_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L2SB_size11_3_sram_inv[0:3]));

	mux_tree_tapbuf_L2SB_size11_mem mem_left_track_29 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size12_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size11_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size11_4_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L2SB_size11_4_sram_inv[0:3]));

	mux_tree_tapbuf_L2SB_size11_mem mem_left_track_33 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size11_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size11_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size11_5_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L2SB_size11_5_sram_inv[0:3]));

	mux_tree_tapbuf_L2SB_size11_mem mem_left_track_37 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size11_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size11_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size11_6_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L2SB_size11_6_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size17 mux_right_track_38 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_8__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_26__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_32__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_34__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_40__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_46__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_52__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_54__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_60__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_66__pin_a2f_o_0_, chany_bottom_in[18], chany_bottom_in[48], chany_bottom_in[78], chanx_left_in[20], chanx_left_in[60]}),
		.sram(mux_tree_tapbuf_L4SB_size17_0_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_L4SB_size17_0_sram_inv[0:4]),
		.out(chanx_right_out[19]));

	mux_tree_tapbuf_L4SB_size17 mux_right_track_46 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_9__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_27__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_33__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_35__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_41__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_47__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_53__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_55__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_61__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_67__pin_a2f_o_0_, chany_bottom_in[17], chany_bottom_in[47], chany_bottom_in[77], chanx_left_in[21], chanx_left_in[61]}),
		.sram(mux_tree_tapbuf_L4SB_size17_1_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_L4SB_size17_1_sram_inv[0:4]),
		.out(chanx_right_out[23]));

	mux_tree_tapbuf_L4SB_size17 mux_right_track_54 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_10__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_28__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_34__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_36__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_42__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_48__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_54__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_56__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_62__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_68__pin_a2f_o_0_, chany_bottom_in[16], chany_bottom_in[46], chany_bottom_in[76], chanx_left_in[23], chanx_left_in[63]}),
		.sram(mux_tree_tapbuf_L4SB_size17_2_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_L4SB_size17_2_sram_inv[0:4]),
		.out(chanx_right_out[27]));

	mux_tree_tapbuf_L4SB_size17 mux_right_track_62 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_11__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_29__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_35__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_37__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_43__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_49__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_55__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_57__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_63__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_69__pin_a2f_o_0_, chany_bottom_in[15], chany_bottom_in[45], chany_bottom_in[75], chanx_left_in[24], chanx_left_in[64]}),
		.sram(mux_tree_tapbuf_L4SB_size17_3_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_L4SB_size17_3_sram_inv[0:4]),
		.out(chanx_right_out[31]));

	mux_tree_tapbuf_L4SB_size17 mux_right_track_70 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_24__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_30__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_36__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_38__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_44__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_50__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_56__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_58__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_64__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_70__pin_a2f_o_0_, chany_bottom_in[14], chany_bottom_in[44], chany_bottom_in[74], chanx_left_in[25], chanx_left_in[65]}),
		.sram(mux_tree_tapbuf_L4SB_size17_4_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_L4SB_size17_4_sram_inv[0:4]),
		.out(chanx_right_out[35]));

	mux_tree_tapbuf_L4SB_size17 mux_right_track_78 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_25__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_31__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_37__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_39__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_45__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_51__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_57__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_59__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_65__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_71__pin_a2f_o_0_, chany_bottom_in[13], chany_bottom_in[43], chany_bottom_in[73], chanx_left_in[27], chanx_left_in[67]}),
		.sram(mux_tree_tapbuf_L4SB_size17_5_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_L4SB_size17_5_sram_inv[0:4]),
		.out(chanx_right_out[39]));

	mux_tree_tapbuf_L4SB_size17 mux_right_track_86 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_8__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_26__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_32__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_38__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_40__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_46__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_52__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_58__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_60__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_66__pin_a2f_o_0_, chany_bottom_in[12], chany_bottom_in[42], chany_bottom_in[72], chanx_left_in[28], chanx_left_in[68]}),
		.sram(mux_tree_tapbuf_L4SB_size17_6_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_L4SB_size17_6_sram_inv[0:4]),
		.out(chanx_right_out[43]));

	mux_tree_tapbuf_L4SB_size17 mux_right_track_94 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_9__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_27__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_33__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_39__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_41__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_47__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_53__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_59__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_61__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_67__pin_a2f_o_0_, chany_bottom_in[11], chany_bottom_in[41], chany_bottom_in[71], chanx_left_in[29], chanx_left_in[69]}),
		.sram(mux_tree_tapbuf_L4SB_size17_7_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_L4SB_size17_7_sram_inv[0:4]),
		.out(chanx_right_out[47]));

	mux_tree_tapbuf_L4SB_size17 mux_right_track_102 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_8__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_10__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_28__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_34__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_40__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_42__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_48__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_54__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_60__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_62__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_68__pin_a2f_o_0_, chany_bottom_in[10], chany_bottom_in[40], chany_bottom_in[70], chanx_left_in[31], chanx_left_in[71]}),
		.sram(mux_tree_tapbuf_L4SB_size17_8_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_L4SB_size17_8_sram_inv[0:4]),
		.out(chanx_right_out[51]));

	mux_tree_tapbuf_L4SB_size17 mux_right_track_110 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_9__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_11__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_29__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_35__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_41__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_43__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_49__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_55__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_61__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_63__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_69__pin_a2f_o_0_, chany_bottom_in[9], chany_bottom_in[39], chany_bottom_in[69], chanx_left_in[32], chanx_left_in[72]}),
		.sram(mux_tree_tapbuf_L4SB_size17_9_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_L4SB_size17_9_sram_inv[0:4]),
		.out(chanx_right_out[55]));

	mux_tree_tapbuf_L4SB_size17 mux_right_track_118 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_10__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_24__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_30__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_36__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_42__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_44__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_50__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_56__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_62__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_64__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_70__pin_a2f_o_0_, chany_bottom_in[8], chany_bottom_in[38], chany_bottom_in[68], chanx_left_in[33], chanx_left_in[73]}),
		.sram(mux_tree_tapbuf_L4SB_size17_10_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_L4SB_size17_10_sram_inv[0:4]),
		.out(chanx_right_out[59]));

	mux_tree_tapbuf_L4SB_size17 mux_right_track_126 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_11__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_25__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_31__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_37__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_43__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_45__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_51__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_57__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_63__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_65__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_71__pin_a2f_o_0_, chany_bottom_in[7], chany_bottom_in[37], chany_bottom_in[67], chanx_left_in[35], chanx_left_in[75]}),
		.sram(mux_tree_tapbuf_L4SB_size17_11_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_L4SB_size17_11_sram_inv[0:4]),
		.out(chanx_right_out[63]));

	mux_tree_tapbuf_L4SB_size17 mux_right_track_134 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_24__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_26__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_32__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_38__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_44__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_46__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_52__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_58__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_64__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_66__pin_a2f_o_0_, chany_bottom_in[6], chany_bottom_in[36], chany_bottom_in[66], chanx_left_in[36], chanx_left_in[76]}),
		.sram(mux_tree_tapbuf_L4SB_size17_12_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_L4SB_size17_12_sram_inv[0:4]),
		.out(chanx_right_out[67]));

	mux_tree_tapbuf_L4SB_size17 mux_right_track_190 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_25__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_31__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_33__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_39__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_45__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_51__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_53__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_59__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_65__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_71__pin_a2f_o_0_, chany_bottom_in[29], chany_bottom_in[59], chany_bottom_in[89], chanx_left_in[45], chanx_left_in[85]}),
		.sram(mux_tree_tapbuf_L4SB_size17_13_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_L4SB_size17_13_sram_inv[0:4]),
		.out(chanx_right_out[95]));

	mux_tree_tapbuf_L4SB_size17 mux_left_track_39 (
		.in({chanx_right_in[20], chanx_right_in[60], chany_bottom_in[9], chany_bottom_in[39], chany_bottom_in[69], left_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_8__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_26__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_32__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_34__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_40__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_46__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_52__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_54__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_60__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_66__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size17_14_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_L4SB_size17_14_sram_inv[0:4]),
		.out(chanx_left_out[19]));

	mux_tree_tapbuf_L4SB_size17 mux_left_track_47 (
		.in({chanx_right_in[21], chanx_right_in[61], chany_bottom_in[10], chany_bottom_in[40], chany_bottom_in[70], left_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_9__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_27__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_33__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_35__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_41__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_47__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_53__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_55__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_61__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_67__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size17_15_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_L4SB_size17_15_sram_inv[0:4]),
		.out(chanx_left_out[23]));

	mux_tree_tapbuf_L4SB_size17 mux_left_track_55 (
		.in({chanx_right_in[23], chanx_right_in[63], chany_bottom_in[11], chany_bottom_in[41], chany_bottom_in[71], left_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_10__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_28__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_34__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_36__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_42__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_48__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_54__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_56__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_62__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_68__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size17_16_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_L4SB_size17_16_sram_inv[0:4]),
		.out(chanx_left_out[27]));

	mux_tree_tapbuf_L4SB_size17 mux_left_track_63 (
		.in({chanx_right_in[24], chanx_right_in[64], chany_bottom_in[12], chany_bottom_in[42], chany_bottom_in[72], left_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_11__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_29__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_35__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_37__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_43__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_49__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_55__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_57__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_63__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_69__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size17_17_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_L4SB_size17_17_sram_inv[0:4]),
		.out(chanx_left_out[31]));

	mux_tree_tapbuf_L4SB_size17 mux_left_track_71 (
		.in({chanx_right_in[25], chanx_right_in[65], chany_bottom_in[13], chany_bottom_in[43], chany_bottom_in[73], left_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_24__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_30__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_36__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_38__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_44__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_50__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_56__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_58__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_64__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_70__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size17_18_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_L4SB_size17_18_sram_inv[0:4]),
		.out(chanx_left_out[35]));

	mux_tree_tapbuf_L4SB_size17 mux_left_track_79 (
		.in({chanx_right_in[27], chanx_right_in[67], chany_bottom_in[14], chany_bottom_in[44], chany_bottom_in[74], left_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_25__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_31__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_37__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_39__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_45__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_51__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_57__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_59__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_65__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_71__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size17_19_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_L4SB_size17_19_sram_inv[0:4]),
		.out(chanx_left_out[39]));

	mux_tree_tapbuf_L4SB_size17 mux_left_track_87 (
		.in({chanx_right_in[28], chanx_right_in[68], chany_bottom_in[15], chany_bottom_in[45], chany_bottom_in[75], left_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_8__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_26__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_32__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_38__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_40__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_46__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_52__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_58__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_60__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_66__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size17_20_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_L4SB_size17_20_sram_inv[0:4]),
		.out(chanx_left_out[43]));

	mux_tree_tapbuf_L4SB_size17 mux_left_track_95 (
		.in({chanx_right_in[29], chanx_right_in[69], chany_bottom_in[16], chany_bottom_in[46], chany_bottom_in[76], left_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_9__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_27__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_33__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_39__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_41__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_47__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_53__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_59__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_61__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_67__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size17_21_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_L4SB_size17_21_sram_inv[0:4]),
		.out(chanx_left_out[47]));

	mux_tree_tapbuf_L4SB_size17 mux_left_track_103 (
		.in({chanx_right_in[31], chanx_right_in[71], chany_bottom_in[17], chany_bottom_in[47], chany_bottom_in[77], left_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_8__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_10__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_28__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_34__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_40__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_42__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_48__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_54__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_60__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_62__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_68__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size17_22_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_L4SB_size17_22_sram_inv[0:4]),
		.out(chanx_left_out[51]));

	mux_tree_tapbuf_L4SB_size17 mux_left_track_111 (
		.in({chanx_right_in[32], chanx_right_in[72], chany_bottom_in[18], chany_bottom_in[48], chany_bottom_in[78], left_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_9__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_11__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_29__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_35__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_41__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_43__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_49__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_55__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_61__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_63__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_69__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size17_23_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_L4SB_size17_23_sram_inv[0:4]),
		.out(chanx_left_out[55]));

	mux_tree_tapbuf_L4SB_size17 mux_left_track_119 (
		.in({chanx_right_in[33], chanx_right_in[73], chany_bottom_in[19], chany_bottom_in[49], chany_bottom_in[79], left_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_10__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_24__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_30__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_36__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_42__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_44__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_50__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_56__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_62__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_64__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_70__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size17_24_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_L4SB_size17_24_sram_inv[0:4]),
		.out(chanx_left_out[59]));

	mux_tree_tapbuf_L4SB_size17 mux_left_track_127 (
		.in({chanx_right_in[35], chanx_right_in[75], chany_bottom_in[20], chany_bottom_in[50], chany_bottom_in[80], left_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_11__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_25__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_31__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_37__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_43__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_45__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_51__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_57__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_63__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_65__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_71__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size17_25_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_L4SB_size17_25_sram_inv[0:4]),
		.out(chanx_left_out[63]));

	mux_tree_tapbuf_L4SB_size17 mux_left_track_135 (
		.in({chanx_right_in[36], chanx_right_in[76], chany_bottom_in[21], chany_bottom_in[51], chany_bottom_in[81], left_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_24__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_26__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_32__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_38__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_44__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_46__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_52__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_58__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_64__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_66__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size17_26_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_L4SB_size17_26_sram_inv[0:4]),
		.out(chanx_left_out[67]));

	mux_tree_tapbuf_L4SB_size17 mux_left_track_143 (
		.in({chanx_right_in[37], chanx_right_in[77], chany_bottom_in[22], chany_bottom_in[52], chany_bottom_in[82], left_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_25__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_27__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_33__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_39__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_45__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_47__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_53__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_59__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_65__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_67__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size17_27_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_L4SB_size17_27_sram_inv[0:4]),
		.out(chanx_left_out[71]));

	mux_tree_tapbuf_L4SB_size17 mux_left_track_151 (
		.in({chanx_right_in[39], chanx_right_in[79], chany_bottom_in[23], chany_bottom_in[53], chany_bottom_in[83], left_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_8__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_26__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_28__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_34__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_40__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_46__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_48__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_54__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_60__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_66__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_68__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size17_28_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_L4SB_size17_28_sram_inv[0:4]),
		.out(chanx_left_out[75]));

	mux_tree_tapbuf_L4SB_size17 mux_left_track_159 (
		.in({chanx_right_in[40], chanx_right_in[80], chany_bottom_in[24], chany_bottom_in[54], chany_bottom_in[84], left_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_9__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_27__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_29__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_35__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_41__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_47__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_49__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_55__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_61__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_67__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_69__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size17_29_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_L4SB_size17_29_sram_inv[0:4]),
		.out(chanx_left_out[79]));

	mux_tree_tapbuf_L4SB_size17 mux_left_track_167 (
		.in({chanx_right_in[41], chanx_right_in[81], chany_bottom_in[25], chany_bottom_in[55], chany_bottom_in[85], left_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_10__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_28__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_30__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_36__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_42__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_48__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_50__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_56__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_62__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_68__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_70__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size17_30_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_L4SB_size17_30_sram_inv[0:4]),
		.out(chanx_left_out[83]));

	mux_tree_tapbuf_L4SB_size17 mux_left_track_175 (
		.in({chanx_right_in[43], chanx_right_in[83], chany_bottom_in[26], chany_bottom_in[56], chany_bottom_in[86], left_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_11__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_29__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_31__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_37__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_43__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_49__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_51__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_57__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_63__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_69__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_71__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size17_31_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_L4SB_size17_31_sram_inv[0:4]),
		.out(chanx_left_out[87]));

	mux_tree_tapbuf_L4SB_size17 mux_left_track_183 (
		.in({chanx_right_in[44], chanx_right_in[84], chany_bottom_in[27], chany_bottom_in[57], chany_bottom_in[87], left_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_24__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_30__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_32__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_38__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_44__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_50__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_52__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_58__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_64__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_70__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size17_32_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_L4SB_size17_32_sram_inv[0:4]),
		.out(chanx_left_out[91]));

	mux_tree_tapbuf_L4SB_size17 mux_left_track_191 (
		.in({chanx_right_in[45], chanx_right_in[85], chany_bottom_in[28], chany_bottom_in[58], chany_bottom_in[88], left_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_25__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_31__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_33__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_39__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_45__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_51__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_53__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_59__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_65__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_71__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size17_33_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_L4SB_size17_33_sram_inv[0:4]),
		.out(chanx_left_out[95]));

	mux_tree_tapbuf_L4SB_size17_mem mem_right_track_38 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size11_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size17_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size17_0_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_L4SB_size17_0_sram_inv[0:4]));

	mux_tree_tapbuf_L4SB_size17_mem mem_right_track_46 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size17_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size17_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size17_1_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_L4SB_size17_1_sram_inv[0:4]));

	mux_tree_tapbuf_L4SB_size17_mem mem_right_track_54 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size17_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size17_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size17_2_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_L4SB_size17_2_sram_inv[0:4]));

	mux_tree_tapbuf_L4SB_size17_mem mem_right_track_62 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size17_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size17_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size17_3_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_L4SB_size17_3_sram_inv[0:4]));

	mux_tree_tapbuf_L4SB_size17_mem mem_right_track_70 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size17_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size17_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size17_4_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_L4SB_size17_4_sram_inv[0:4]));

	mux_tree_tapbuf_L4SB_size17_mem mem_right_track_78 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size17_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size17_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size17_5_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_L4SB_size17_5_sram_inv[0:4]));

	mux_tree_tapbuf_L4SB_size17_mem mem_right_track_86 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size17_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size17_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size17_6_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_L4SB_size17_6_sram_inv[0:4]));

	mux_tree_tapbuf_L4SB_size17_mem mem_right_track_94 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size17_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size17_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size17_7_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_L4SB_size17_7_sram_inv[0:4]));

	mux_tree_tapbuf_L4SB_size17_mem mem_right_track_102 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size17_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size17_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size17_8_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_L4SB_size17_8_sram_inv[0:4]));

	mux_tree_tapbuf_L4SB_size17_mem mem_right_track_110 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size17_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size17_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size17_9_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_L4SB_size17_9_sram_inv[0:4]));

	mux_tree_tapbuf_L4SB_size17_mem mem_right_track_118 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size17_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size17_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size17_10_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_L4SB_size17_10_sram_inv[0:4]));

	mux_tree_tapbuf_L4SB_size17_mem mem_right_track_126 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size17_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size17_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size17_11_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_L4SB_size17_11_sram_inv[0:4]));

	mux_tree_tapbuf_L4SB_size17_mem mem_right_track_134 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size17_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size17_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size17_12_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_L4SB_size17_12_sram_inv[0:4]));

	mux_tree_tapbuf_L4SB_size17_mem mem_right_track_190 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size18_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size17_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size17_13_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_L4SB_size17_13_sram_inv[0:4]));

	mux_tree_tapbuf_L4SB_size17_mem mem_left_track_39 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size11_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size17_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size17_14_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_L4SB_size17_14_sram_inv[0:4]));

	mux_tree_tapbuf_L4SB_size17_mem mem_left_track_47 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size17_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size17_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size17_15_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_L4SB_size17_15_sram_inv[0:4]));

	mux_tree_tapbuf_L4SB_size17_mem mem_left_track_55 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size17_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size17_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size17_16_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_L4SB_size17_16_sram_inv[0:4]));

	mux_tree_tapbuf_L4SB_size17_mem mem_left_track_63 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size17_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size17_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size17_17_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_L4SB_size17_17_sram_inv[0:4]));

	mux_tree_tapbuf_L4SB_size17_mem mem_left_track_71 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size17_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size17_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size17_18_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_L4SB_size17_18_sram_inv[0:4]));

	mux_tree_tapbuf_L4SB_size17_mem mem_left_track_79 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size17_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size17_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size17_19_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_L4SB_size17_19_sram_inv[0:4]));

	mux_tree_tapbuf_L4SB_size17_mem mem_left_track_87 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size17_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size17_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size17_20_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_L4SB_size17_20_sram_inv[0:4]));

	mux_tree_tapbuf_L4SB_size17_mem mem_left_track_95 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size17_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size17_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size17_21_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_L4SB_size17_21_sram_inv[0:4]));

	mux_tree_tapbuf_L4SB_size17_mem mem_left_track_103 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size17_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size17_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size17_22_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_L4SB_size17_22_sram_inv[0:4]));

	mux_tree_tapbuf_L4SB_size17_mem mem_left_track_111 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size17_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size17_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size17_23_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_L4SB_size17_23_sram_inv[0:4]));

	mux_tree_tapbuf_L4SB_size17_mem mem_left_track_119 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size17_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size17_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size17_24_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_L4SB_size17_24_sram_inv[0:4]));

	mux_tree_tapbuf_L4SB_size17_mem mem_left_track_127 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size17_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size17_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size17_25_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_L4SB_size17_25_sram_inv[0:4]));

	mux_tree_tapbuf_L4SB_size17_mem mem_left_track_135 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size17_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size17_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size17_26_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_L4SB_size17_26_sram_inv[0:4]));

	mux_tree_tapbuf_L4SB_size17_mem mem_left_track_143 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size17_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size17_mem_27_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size17_27_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_L4SB_size17_27_sram_inv[0:4]));

	mux_tree_tapbuf_L4SB_size17_mem mem_left_track_151 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size17_mem_27_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size17_mem_28_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size17_28_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_L4SB_size17_28_sram_inv[0:4]));

	mux_tree_tapbuf_L4SB_size17_mem mem_left_track_159 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size17_mem_28_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size17_mem_29_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size17_29_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_L4SB_size17_29_sram_inv[0:4]));

	mux_tree_tapbuf_L4SB_size17_mem mem_left_track_167 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size17_mem_29_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size17_mem_30_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size17_30_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_L4SB_size17_30_sram_inv[0:4]));

	mux_tree_tapbuf_L4SB_size17_mem mem_left_track_175 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size17_mem_30_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size17_mem_31_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size17_31_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_L4SB_size17_31_sram_inv[0:4]));

	mux_tree_tapbuf_L4SB_size17_mem mem_left_track_183 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size17_mem_31_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size17_mem_32_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size17_32_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_L4SB_size17_32_sram_inv[0:4]));

	mux_tree_tapbuf_L4SB_size17_mem mem_left_track_191 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size17_mem_32_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size17_33_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_L4SB_size17_33_sram_inv[0:4]));

	mux_tree_tapbuf_L4SB_size18 mux_right_track_142 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_25__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_27__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_33__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_39__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_45__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_47__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_53__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_59__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_65__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_67__pin_a2f_o_0_, chany_bottom_in[5], chany_bottom_in[35], chany_bottom_in[65], chany_bottom_in[95], chanx_left_in[37], chanx_left_in[77]}),
		.sram(mux_tree_tapbuf_L4SB_size18_0_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_L4SB_size18_0_sram_inv[0:4]),
		.out(chanx_right_out[71]));

	mux_tree_tapbuf_L4SB_size18 mux_right_track_150 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_8__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_26__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_28__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_34__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_40__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_46__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_48__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_54__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_60__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_66__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_68__pin_a2f_o_0_, chany_bottom_in[4], chany_bottom_in[34], chany_bottom_in[64], chany_bottom_in[94], chanx_left_in[39], chanx_left_in[79]}),
		.sram(mux_tree_tapbuf_L4SB_size18_1_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_L4SB_size18_1_sram_inv[0:4]),
		.out(chanx_right_out[75]));

	mux_tree_tapbuf_L4SB_size18 mux_right_track_158 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_9__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_27__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_29__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_35__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_41__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_47__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_49__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_55__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_61__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_67__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_69__pin_a2f_o_0_, chany_bottom_in[3], chany_bottom_in[33], chany_bottom_in[63], chany_bottom_in[93], chanx_left_in[40], chanx_left_in[80]}),
		.sram(mux_tree_tapbuf_L4SB_size18_2_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_L4SB_size18_2_sram_inv[0:4]),
		.out(chanx_right_out[79]));

	mux_tree_tapbuf_L4SB_size18 mux_right_track_166 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_10__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_28__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_30__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_36__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_42__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_48__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_50__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_56__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_62__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_68__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_70__pin_a2f_o_0_, chany_bottom_in[2], chany_bottom_in[32], chany_bottom_in[62], chany_bottom_in[92], chanx_left_in[41], chanx_left_in[81]}),
		.sram(mux_tree_tapbuf_L4SB_size18_3_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_L4SB_size18_3_sram_inv[0:4]),
		.out(chanx_right_out[83]));

	mux_tree_tapbuf_L4SB_size18 mux_right_track_174 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_11__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_29__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_31__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_37__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_43__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_49__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_51__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_57__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_63__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_69__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_71__pin_a2f_o_0_, chany_bottom_in[1], chany_bottom_in[31], chany_bottom_in[61], chany_bottom_in[91], chanx_left_in[43], chanx_left_in[83]}),
		.sram(mux_tree_tapbuf_L4SB_size18_4_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_L4SB_size18_4_sram_inv[0:4]),
		.out(chanx_right_out[87]));

	mux_tree_tapbuf_L4SB_size18 mux_right_track_182 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_24__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_30__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_32__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_38__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_44__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_50__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_52__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_58__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_64__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_70__pin_a2f_o_0_, chany_bottom_in[0], chany_bottom_in[30], chany_bottom_in[60], chany_bottom_in[90], chanx_left_in[44], chanx_left_in[84]}),
		.sram(mux_tree_tapbuf_L4SB_size18_5_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_L4SB_size18_5_sram_inv[0:4]),
		.out(chanx_right_out[91]));

	mux_tree_tapbuf_L4SB_size18_mem mem_right_track_142 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size17_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size18_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size18_0_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_L4SB_size18_0_sram_inv[0:4]));

	mux_tree_tapbuf_L4SB_size18_mem mem_right_track_150 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size18_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size18_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size18_1_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_L4SB_size18_1_sram_inv[0:4]));

	mux_tree_tapbuf_L4SB_size18_mem mem_right_track_158 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size18_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size18_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size18_2_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_L4SB_size18_2_sram_inv[0:4]));

	mux_tree_tapbuf_L4SB_size18_mem mem_right_track_166 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size18_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size18_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size18_3_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_L4SB_size18_3_sram_inv[0:4]));

	mux_tree_tapbuf_L4SB_size18_mem mem_right_track_174 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size18_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size18_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size18_4_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_L4SB_size18_4_sram_inv[0:4]));

	mux_tree_tapbuf_L4SB_size18_mem mem_right_track_182 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size18_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size18_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size18_5_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_L4SB_size18_5_sram_inv[0:4]));

	mux_tree_tapbuf_L2SB_size4 mux_bottom_track_1 (
		.in({chanx_right_in[0], bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_, chanx_left_in[0], chanx_left_in[3]}),
		.sram(mux_tree_tapbuf_L2SB_size4_0_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_0_sram_inv[0:1]),
		.out(chany_bottom_out[0]));

	mux_tree_tapbuf_L2SB_size4 mux_bottom_track_3 (
		.in({chanx_right_in[2], bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_, chanx_left_in[2], chanx_left_in[5]}),
		.sram(mux_tree_tapbuf_L2SB_size4_1_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_1_sram_inv[0:1]),
		.out(chany_bottom_out[1]));

	mux_tree_tapbuf_L2SB_size4 mux_bottom_track_5 (
		.in({chanx_right_in[4], bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_, chanx_left_in[4], chanx_left_in[7]}),
		.sram(mux_tree_tapbuf_L2SB_size4_2_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_2_sram_inv[0:1]),
		.out(chany_bottom_out[2]));

	mux_tree_tapbuf_L2SB_size4 mux_bottom_track_7 (
		.in({chanx_right_in[6], bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_, chanx_left_in[6], chanx_left_in[9]}),
		.sram(mux_tree_tapbuf_L2SB_size4_3_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_3_sram_inv[0:1]),
		.out(chany_bottom_out[3]));

	mux_tree_tapbuf_L2SB_size4 mux_bottom_track_9 (
		.in({chanx_right_in[8], bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_, chanx_left_in[8], chanx_left_in[11]}),
		.sram(mux_tree_tapbuf_L2SB_size4_4_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_4_sram_inv[0:1]),
		.out(chany_bottom_out[4]));

	mux_tree_tapbuf_L2SB_size4 mux_bottom_track_11 (
		.in({chanx_right_in[10], bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_, chanx_left_in[10], chanx_left_in[13]}),
		.sram(mux_tree_tapbuf_L2SB_size4_5_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_5_sram_inv[0:1]),
		.out(chany_bottom_out[5]));

	mux_tree_tapbuf_L2SB_size4 mux_bottom_track_13 (
		.in({chanx_right_in[12], bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_, chanx_left_in[12], chanx_left_in[15]}),
		.sram(mux_tree_tapbuf_L2SB_size4_6_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_6_sram_inv[0:1]),
		.out(chany_bottom_out[6]));

	mux_tree_tapbuf_L2SB_size4 mux_bottom_track_15 (
		.in({chanx_right_in[14], bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_, chanx_left_in[14], chanx_left_in[17]}),
		.sram(mux_tree_tapbuf_L2SB_size4_7_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_7_sram_inv[0:1]),
		.out(chany_bottom_out[7]));

	mux_tree_tapbuf_L2SB_size4 mux_bottom_track_17 (
		.in({chanx_right_in[16], bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_, chanx_left_in[16], chanx_left_in[18]}),
		.sram(mux_tree_tapbuf_L2SB_size4_8_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_8_sram_inv[0:1]),
		.out(chany_bottom_out[8]));

	mux_tree_tapbuf_L2SB_size4 mux_bottom_track_19 (
		.in({chanx_right_in[19], bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_, chanx_left_in[19], chanx_left_in[22]}),
		.sram(mux_tree_tapbuf_L2SB_size4_9_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_9_sram_inv[0:1]),
		.out(chany_bottom_out[9]));

	mux_tree_tapbuf_L2SB_size4 mux_bottom_track_21 (
		.in({chanx_right_in[20], bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_, chanx_left_in[20], chanx_left_in[26]}),
		.sram(mux_tree_tapbuf_L2SB_size4_10_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_10_sram_inv[0:1]),
		.out(chany_bottom_out[10]));

	mux_tree_tapbuf_L2SB_size4 mux_bottom_track_23 (
		.in({chanx_right_in[21], bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_, chanx_left_in[21], chanx_left_in[30]}),
		.sram(mux_tree_tapbuf_L2SB_size4_11_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_11_sram_inv[0:1]),
		.out(chany_bottom_out[11]));

	mux_tree_tapbuf_L2SB_size4_mem mem_bottom_track_1 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size17_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_0_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_0_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_bottom_track_3 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_1_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_1_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_bottom_track_5 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_2_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_2_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_bottom_track_7 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_3_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_3_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_bottom_track_9 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_4_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_4_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_bottom_track_11 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_5_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_5_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_bottom_track_13 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_6_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_6_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_bottom_track_15 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_7_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_7_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_bottom_track_17 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_8_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_8_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_bottom_track_19 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_9_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_9_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_bottom_track_21 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_10_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_10_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_bottom_track_23 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_11_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_11_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size3 mux_bottom_track_25 (
		.in({chanx_right_in[23], chanx_left_in[23], chanx_left_in[34]}),
		.sram(mux_tree_tapbuf_L2SB_size3_0_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size3_0_sram_inv[0:1]),
		.out(chany_bottom_out[12]));

	mux_tree_tapbuf_L2SB_size3 mux_bottom_track_27 (
		.in({chanx_right_in[24], chanx_left_in[24], chanx_left_in[38]}),
		.sram(mux_tree_tapbuf_L2SB_size3_1_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size3_1_sram_inv[0:1]),
		.out(chany_bottom_out[13]));

	mux_tree_tapbuf_L2SB_size3 mux_bottom_track_29 (
		.in({chanx_right_in[25], chanx_left_in[25], chanx_left_in[42]}),
		.sram(mux_tree_tapbuf_L2SB_size3_2_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size3_2_sram_inv[0:1]),
		.out(chany_bottom_out[14]));

	mux_tree_tapbuf_L2SB_size3 mux_bottom_track_31 (
		.in({chanx_right_in[27], chanx_left_in[27], chanx_left_in[46]}),
		.sram(mux_tree_tapbuf_L2SB_size3_3_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size3_3_sram_inv[0:1]),
		.out(chany_bottom_out[15]));

	mux_tree_tapbuf_L2SB_size3 mux_bottom_track_33 (
		.in({chanx_right_in[28], chanx_left_in[28], chanx_left_in[50]}),
		.sram(mux_tree_tapbuf_L2SB_size3_4_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size3_4_sram_inv[0:1]),
		.out(chany_bottom_out[16]));

	mux_tree_tapbuf_L2SB_size3 mux_bottom_track_35 (
		.in({chanx_right_in[29], chanx_left_in[29], chanx_left_in[54]}),
		.sram(mux_tree_tapbuf_L2SB_size3_5_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size3_5_sram_inv[0:1]),
		.out(chany_bottom_out[17]));

	mux_tree_tapbuf_L2SB_size3 mux_bottom_track_37 (
		.in({chanx_right_in[31], chanx_left_in[31], chanx_left_in[58]}),
		.sram(mux_tree_tapbuf_L2SB_size3_6_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size3_6_sram_inv[0:1]),
		.out(chany_bottom_out[18]));

	mux_tree_tapbuf_L2SB_size3_mem mem_bottom_track_25 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size3_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size3_0_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size3_0_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size3_mem mem_bottom_track_27 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size3_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size3_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size3_1_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size3_1_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size3_mem mem_bottom_track_29 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size3_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size3_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size3_2_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size3_2_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size3_mem mem_bottom_track_31 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size3_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size3_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size3_3_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size3_3_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size3_mem mem_bottom_track_33 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size3_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size3_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size3_4_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size3_4_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size3_mem mem_bottom_track_35 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size3_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size3_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size3_5_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size3_5_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size3_mem mem_bottom_track_37 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size3_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size3_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size3_6_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size3_6_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size5 mux_bottom_track_39 (
		.in({chanx_right_in[32], bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_, chanx_left_in[32], chanx_left_in[62]}),
		.sram(mux_tree_tapbuf_L4SB_size5_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_0_sram_inv[0:2]),
		.out(chany_bottom_out[19]));

	mux_tree_tapbuf_L4SB_size5 mux_bottom_track_41 (
		.in({chanx_right_in[33], bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_, chanx_left_in[33], chanx_left_in[66]}),
		.sram(mux_tree_tapbuf_L4SB_size5_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_1_sram_inv[0:2]),
		.out(chany_bottom_out[20]));

	mux_tree_tapbuf_L4SB_size5 mux_bottom_track_43 (
		.in({chanx_right_in[35], bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_, chanx_left_in[35], chanx_left_in[70]}),
		.sram(mux_tree_tapbuf_L4SB_size5_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_2_sram_inv[0:2]),
		.out(chany_bottom_out[21]));

	mux_tree_tapbuf_L4SB_size5 mux_bottom_track_45 (
		.in({chanx_right_in[36], bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_, chanx_left_in[36], chanx_left_in[74]}),
		.sram(mux_tree_tapbuf_L4SB_size5_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_3_sram_inv[0:2]),
		.out(chany_bottom_out[22]));

	mux_tree_tapbuf_L4SB_size5 mux_bottom_track_47 (
		.in({chanx_right_in[37], bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_, chanx_left_in[37], chanx_left_in[78]}),
		.sram(mux_tree_tapbuf_L4SB_size5_4_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_4_sram_inv[0:2]),
		.out(chany_bottom_out[23]));

	mux_tree_tapbuf_L4SB_size5 mux_bottom_track_53 (
		.in({chanx_right_in[41], bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_, chanx_left_in[41], chanx_left_in[90]}),
		.sram(mux_tree_tapbuf_L4SB_size5_5_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_5_sram_inv[0:2]),
		.out(chany_bottom_out[26]));

	mux_tree_tapbuf_L4SB_size5 mux_bottom_track_55 (
		.in({chanx_right_in[43], bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_, chanx_left_in[43], chanx_left_in[94]}),
		.sram(mux_tree_tapbuf_L4SB_size5_6_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_6_sram_inv[0:2]),
		.out(chany_bottom_out[27]));

	mux_tree_tapbuf_L4SB_size5 mux_bottom_track_57 (
		.in({chanx_right_in[44], bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_, chanx_left_in[44], chanx_left_in[95]}),
		.sram(mux_tree_tapbuf_L4SB_size5_7_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_7_sram_inv[0:2]),
		.out(chany_bottom_out[28]));

	mux_tree_tapbuf_L4SB_size5 mux_bottom_track_131 (
		.in({chanx_right_in[93], chanx_right_in[95], bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_, chanx_left_in[93]}),
		.sram(mux_tree_tapbuf_L4SB_size5_8_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_8_sram_inv[0:2]),
		.out(chany_bottom_out[65]));

	mux_tree_tapbuf_L4SB_size5_mem mem_bottom_track_39 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size3_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size5_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size5_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_0_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size5_mem mem_bottom_track_41 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size5_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size5_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size5_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_1_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size5_mem mem_bottom_track_43 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size5_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size5_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size5_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_2_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size5_mem mem_bottom_track_45 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size5_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size5_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size5_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_3_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size5_mem mem_bottom_track_47 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size5_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size5_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size5_4_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_4_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size5_mem mem_bottom_track_53 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size4_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size5_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size5_5_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_5_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size5_mem mem_bottom_track_55 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size5_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size5_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size5_6_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_6_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size5_mem mem_bottom_track_57 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size5_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size5_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size5_7_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_7_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size5_mem mem_bottom_track_131 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size4_mem_27_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size5_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size5_8_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_8_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size4 mux_bottom_track_49 (
		.in({chanx_right_in[39], bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_, chanx_left_in[39], chanx_left_in[82]}),
		.sram(mux_tree_tapbuf_L4SB_size4_0_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_0_sram_inv[0:1]),
		.out(chany_bottom_out[24]));

	mux_tree_tapbuf_L4SB_size4 mux_bottom_track_51 (
		.in({chanx_right_in[40], bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_, chanx_left_in[40], chanx_left_in[86]}),
		.sram(mux_tree_tapbuf_L4SB_size4_1_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_1_sram_inv[0:1]),
		.out(chany_bottom_out[25]));

	mux_tree_tapbuf_L4SB_size4 mux_bottom_track_59 (
		.in({chanx_right_in[45], bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_, chanx_left_in[45]}),
		.sram(mux_tree_tapbuf_L4SB_size4_2_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_2_sram_inv[0:1]),
		.out(chany_bottom_out[29]));

	mux_tree_tapbuf_L4SB_size4 mux_bottom_track_61 (
		.in({chanx_right_in[47], bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_, chanx_left_in[47]}),
		.sram(mux_tree_tapbuf_L4SB_size4_3_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_3_sram_inv[0:1]),
		.out(chany_bottom_out[30]));

	mux_tree_tapbuf_L4SB_size4 mux_bottom_track_67 (
		.in({chanx_right_in[51], bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_, chanx_left_in[51]}),
		.sram(mux_tree_tapbuf_L4SB_size4_4_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_4_sram_inv[0:1]),
		.out(chany_bottom_out[33]));

	mux_tree_tapbuf_L4SB_size4 mux_bottom_track_69 (
		.in({chanx_right_in[52], bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_, chanx_left_in[52]}),
		.sram(mux_tree_tapbuf_L4SB_size4_5_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_5_sram_inv[0:1]),
		.out(chany_bottom_out[34]));

	mux_tree_tapbuf_L4SB_size4 mux_bottom_track_71 (
		.in({chanx_right_in[53], bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_, chanx_left_in[53]}),
		.sram(mux_tree_tapbuf_L4SB_size4_6_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_6_sram_inv[0:1]),
		.out(chany_bottom_out[35]));

	mux_tree_tapbuf_L4SB_size4 mux_bottom_track_73 (
		.in({chanx_right_in[55], bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_, chanx_left_in[55]}),
		.sram(mux_tree_tapbuf_L4SB_size4_7_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_7_sram_inv[0:1]),
		.out(chany_bottom_out[36]));

	mux_tree_tapbuf_L4SB_size4 mux_bottom_track_75 (
		.in({chanx_right_in[56], bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_, chanx_left_in[56]}),
		.sram(mux_tree_tapbuf_L4SB_size4_8_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_8_sram_inv[0:1]),
		.out(chany_bottom_out[37]));

	mux_tree_tapbuf_L4SB_size4 mux_bottom_track_81 (
		.in({chanx_right_in[60], bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_, chanx_left_in[60]}),
		.sram(mux_tree_tapbuf_L4SB_size4_9_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_9_sram_inv[0:1]),
		.out(chany_bottom_out[40]));

	mux_tree_tapbuf_L4SB_size4 mux_bottom_track_83 (
		.in({chanx_right_in[61], bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_, chanx_left_in[61]}),
		.sram(mux_tree_tapbuf_L4SB_size4_10_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_10_sram_inv[0:1]),
		.out(chany_bottom_out[41]));

	mux_tree_tapbuf_L4SB_size4 mux_bottom_track_85 (
		.in({chanx_right_in[63], bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_, chanx_left_in[63]}),
		.sram(mux_tree_tapbuf_L4SB_size4_11_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_11_sram_inv[0:1]),
		.out(chany_bottom_out[42]));

	mux_tree_tapbuf_L4SB_size4 mux_bottom_track_87 (
		.in({chanx_right_in[64], bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_, chanx_left_in[64]}),
		.sram(mux_tree_tapbuf_L4SB_size4_12_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_12_sram_inv[0:1]),
		.out(chany_bottom_out[43]));

	mux_tree_tapbuf_L4SB_size4 mux_bottom_track_89 (
		.in({chanx_right_in[65], bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_, chanx_left_in[65]}),
		.sram(mux_tree_tapbuf_L4SB_size4_13_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_13_sram_inv[0:1]),
		.out(chany_bottom_out[44]));

	mux_tree_tapbuf_L4SB_size4 mux_bottom_track_95 (
		.in({chanx_right_in[69], bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_, chanx_left_in[69]}),
		.sram(mux_tree_tapbuf_L4SB_size4_14_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_14_sram_inv[0:1]),
		.out(chany_bottom_out[47]));

	mux_tree_tapbuf_L4SB_size4 mux_bottom_track_97 (
		.in({chanx_right_in[71], bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_, chanx_left_in[71]}),
		.sram(mux_tree_tapbuf_L4SB_size4_15_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_15_sram_inv[0:1]),
		.out(chany_bottom_out[48]));

	mux_tree_tapbuf_L4SB_size4 mux_bottom_track_99 (
		.in({chanx_right_in[72], bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_, chanx_left_in[72]}),
		.sram(mux_tree_tapbuf_L4SB_size4_16_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_16_sram_inv[0:1]),
		.out(chany_bottom_out[49]));

	mux_tree_tapbuf_L4SB_size4 mux_bottom_track_101 (
		.in({chanx_right_in[73], bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_, chanx_left_in[73]}),
		.sram(mux_tree_tapbuf_L4SB_size4_17_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_17_sram_inv[0:1]),
		.out(chany_bottom_out[50]));

	mux_tree_tapbuf_L4SB_size4 mux_bottom_track_103 (
		.in({chanx_right_in[75], bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_, chanx_left_in[75]}),
		.sram(mux_tree_tapbuf_L4SB_size4_18_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_18_sram_inv[0:1]),
		.out(chany_bottom_out[51]));

	mux_tree_tapbuf_L4SB_size4 mux_bottom_track_109 (
		.in({chanx_right_in[79], bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_, chanx_left_in[79]}),
		.sram(mux_tree_tapbuf_L4SB_size4_19_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_19_sram_inv[0:1]),
		.out(chany_bottom_out[54]));

	mux_tree_tapbuf_L4SB_size4 mux_bottom_track_111 (
		.in({chanx_right_in[80], bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_, chanx_left_in[80]}),
		.sram(mux_tree_tapbuf_L4SB_size4_20_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_20_sram_inv[0:1]),
		.out(chany_bottom_out[55]));

	mux_tree_tapbuf_L4SB_size4 mux_bottom_track_113 (
		.in({chanx_right_in[81], bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_, chanx_left_in[81]}),
		.sram(mux_tree_tapbuf_L4SB_size4_21_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_21_sram_inv[0:1]),
		.out(chany_bottom_out[56]));

	mux_tree_tapbuf_L4SB_size4 mux_bottom_track_115 (
		.in({chanx_right_in[83], bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_, chanx_left_in[83]}),
		.sram(mux_tree_tapbuf_L4SB_size4_22_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_22_sram_inv[0:1]),
		.out(chany_bottom_out[57]));

	mux_tree_tapbuf_L4SB_size4 mux_bottom_track_117 (
		.in({chanx_right_in[84], bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_, chanx_left_in[84]}),
		.sram(mux_tree_tapbuf_L4SB_size4_23_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_23_sram_inv[0:1]),
		.out(chany_bottom_out[58]));

	mux_tree_tapbuf_L4SB_size4 mux_bottom_track_123 (
		.in({chanx_right_in[88], bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_, chanx_left_in[88]}),
		.sram(mux_tree_tapbuf_L4SB_size4_24_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_24_sram_inv[0:1]),
		.out(chany_bottom_out[61]));

	mux_tree_tapbuf_L4SB_size4 mux_bottom_track_125 (
		.in({chanx_right_in[89], bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_, chanx_left_in[89]}),
		.sram(mux_tree_tapbuf_L4SB_size4_25_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_25_sram_inv[0:1]),
		.out(chany_bottom_out[62]));

	mux_tree_tapbuf_L4SB_size4 mux_bottom_track_127 (
		.in({chanx_right_in[91], bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_, chanx_left_in[91]}),
		.sram(mux_tree_tapbuf_L4SB_size4_26_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_26_sram_inv[0:1]),
		.out(chany_bottom_out[63]));

	mux_tree_tapbuf_L4SB_size4 mux_bottom_track_129 (
		.in({chanx_right_in[92], bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_, chanx_left_in[92]}),
		.sram(mux_tree_tapbuf_L4SB_size4_27_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_27_sram_inv[0:1]),
		.out(chany_bottom_out[64]));

	mux_tree_tapbuf_L4SB_size4_mem mem_bottom_track_49 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size5_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size4_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size4_0_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_0_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_bottom_track_51 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size4_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size4_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size4_1_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_1_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_bottom_track_59 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size5_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size4_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size4_2_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_2_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_bottom_track_61 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size4_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size4_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size4_3_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_3_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_bottom_track_67 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size4_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size4_4_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_4_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_bottom_track_69 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size4_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size4_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size4_5_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_5_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_bottom_track_71 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size4_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size4_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size4_6_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_6_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_bottom_track_73 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size4_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size4_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size4_7_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_7_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_bottom_track_75 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size4_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size4_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size4_8_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_8_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_bottom_track_81 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size4_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size4_9_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_9_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_bottom_track_83 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size4_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size4_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size4_10_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_10_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_bottom_track_85 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size4_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size4_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size4_11_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_11_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_bottom_track_87 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size4_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size4_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size4_12_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_12_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_bottom_track_89 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size4_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size4_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size4_13_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_13_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_bottom_track_95 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size4_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size4_14_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_14_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_bottom_track_97 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size4_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size4_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size4_15_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_15_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_bottom_track_99 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size4_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size4_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size4_16_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_16_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_bottom_track_101 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size4_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size4_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size4_17_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_17_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_bottom_track_103 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size4_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size4_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size4_18_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_18_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_bottom_track_109 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size4_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size4_19_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_19_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_bottom_track_111 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size4_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size4_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size4_20_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_20_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_bottom_track_113 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size4_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size4_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size4_21_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_21_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_bottom_track_115 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size4_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size4_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size4_22_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_22_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_bottom_track_117 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size4_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size4_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size4_23_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_23_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_bottom_track_123 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size4_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size4_24_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_24_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_bottom_track_125 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size4_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size4_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size4_25_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_25_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_bottom_track_127 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size4_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size4_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size4_26_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_26_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_bottom_track_129 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size4_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size4_mem_27_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size4_27_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_27_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3 mux_bottom_track_63 (
		.in({chanx_right_in[48], bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_, chanx_left_in[48]}),
		.sram(mux_tree_tapbuf_L4SB_size3_0_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_0_sram_inv[0:1]),
		.out(chany_bottom_out[31]));

	mux_tree_tapbuf_L4SB_size3 mux_bottom_track_65 (
		.in({chanx_right_in[49], bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_, chanx_left_in[49]}),
		.sram(mux_tree_tapbuf_L4SB_size3_1_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_1_sram_inv[0:1]),
		.out(chany_bottom_out[32]));

	mux_tree_tapbuf_L4SB_size3 mux_bottom_track_77 (
		.in({chanx_right_in[57], bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_, chanx_left_in[57]}),
		.sram(mux_tree_tapbuf_L4SB_size3_2_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_2_sram_inv[0:1]),
		.out(chany_bottom_out[38]));

	mux_tree_tapbuf_L4SB_size3 mux_bottom_track_79 (
		.in({chanx_right_in[59], bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_, chanx_left_in[59]}),
		.sram(mux_tree_tapbuf_L4SB_size3_3_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_3_sram_inv[0:1]),
		.out(chany_bottom_out[39]));

	mux_tree_tapbuf_L4SB_size3 mux_bottom_track_91 (
		.in({chanx_right_in[67], bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_, chanx_left_in[67]}),
		.sram(mux_tree_tapbuf_L4SB_size3_4_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_4_sram_inv[0:1]),
		.out(chany_bottom_out[45]));

	mux_tree_tapbuf_L4SB_size3 mux_bottom_track_93 (
		.in({chanx_right_in[68], bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_, chanx_left_in[68]}),
		.sram(mux_tree_tapbuf_L4SB_size3_5_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_5_sram_inv[0:1]),
		.out(chany_bottom_out[46]));

	mux_tree_tapbuf_L4SB_size3 mux_bottom_track_105 (
		.in({chanx_right_in[76], bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_, chanx_left_in[76]}),
		.sram(mux_tree_tapbuf_L4SB_size3_6_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_6_sram_inv[0:1]),
		.out(chany_bottom_out[52]));

	mux_tree_tapbuf_L4SB_size3 mux_bottom_track_107 (
		.in({chanx_right_in[77], bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_, chanx_left_in[77]}),
		.sram(mux_tree_tapbuf_L4SB_size3_7_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_7_sram_inv[0:1]),
		.out(chany_bottom_out[53]));

	mux_tree_tapbuf_L4SB_size3 mux_bottom_track_119 (
		.in({chanx_right_in[85], bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_, chanx_left_in[85]}),
		.sram(mux_tree_tapbuf_L4SB_size3_8_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_8_sram_inv[0:1]),
		.out(chany_bottom_out[59]));

	mux_tree_tapbuf_L4SB_size3 mux_bottom_track_121 (
		.in({chanx_right_in[87], bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_, chanx_left_in[87]}),
		.sram(mux_tree_tapbuf_L4SB_size3_9_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_9_sram_inv[0:1]),
		.out(chany_bottom_out[60]));

	mux_tree_tapbuf_L4SB_size3 mux_bottom_track_137 (
		.in({chanx_right_in[86], bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_10_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_10_sram_inv[0:1]),
		.out(chany_bottom_out[68]));

	mux_tree_tapbuf_L4SB_size3 mux_bottom_track_139 (
		.in({chanx_right_in[82], bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_11_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_11_sram_inv[0:1]),
		.out(chany_bottom_out[69]));

	mux_tree_tapbuf_L4SB_size3 mux_bottom_track_141 (
		.in({chanx_right_in[78], bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_12_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_12_sram_inv[0:1]),
		.out(chany_bottom_out[70]));

	mux_tree_tapbuf_L4SB_size3 mux_bottom_track_143 (
		.in({chanx_right_in[74], bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_13_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_13_sram_inv[0:1]),
		.out(chany_bottom_out[71]));

	mux_tree_tapbuf_L4SB_size3 mux_bottom_track_145 (
		.in({chanx_right_in[70], bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_14_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_14_sram_inv[0:1]),
		.out(chany_bottom_out[72]));

	mux_tree_tapbuf_L4SB_size3 mux_bottom_track_151 (
		.in({chanx_right_in[58], bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_15_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_15_sram_inv[0:1]),
		.out(chany_bottom_out[75]));

	mux_tree_tapbuf_L4SB_size3 mux_bottom_track_153 (
		.in({chanx_right_in[54], bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_16_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_16_sram_inv[0:1]),
		.out(chany_bottom_out[76]));

	mux_tree_tapbuf_L4SB_size3 mux_bottom_track_155 (
		.in({chanx_right_in[50], bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_17_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_17_sram_inv[0:1]),
		.out(chany_bottom_out[77]));

	mux_tree_tapbuf_L4SB_size3 mux_bottom_track_157 (
		.in({chanx_right_in[46], bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_18_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_18_sram_inv[0:1]),
		.out(chany_bottom_out[78]));

	mux_tree_tapbuf_L4SB_size3 mux_bottom_track_159 (
		.in({chanx_right_in[42], bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_19_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_19_sram_inv[0:1]),
		.out(chany_bottom_out[79]));

	mux_tree_tapbuf_L4SB_size3 mux_bottom_track_165 (
		.in({chanx_right_in[30], bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_20_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_20_sram_inv[0:1]),
		.out(chany_bottom_out[82]));

	mux_tree_tapbuf_L4SB_size3 mux_bottom_track_167 (
		.in({chanx_right_in[26], bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_21_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_21_sram_inv[0:1]),
		.out(chany_bottom_out[83]));

	mux_tree_tapbuf_L4SB_size3 mux_bottom_track_169 (
		.in({chanx_right_in[22], bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_22_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_22_sram_inv[0:1]),
		.out(chany_bottom_out[84]));

	mux_tree_tapbuf_L4SB_size3 mux_bottom_track_171 (
		.in({chanx_right_in[18], bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_23_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_23_sram_inv[0:1]),
		.out(chany_bottom_out[85]));

	mux_tree_tapbuf_L4SB_size3 mux_bottom_track_173 (
		.in({chanx_right_in[17], bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_24_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_24_sram_inv[0:1]),
		.out(chany_bottom_out[86]));

	mux_tree_tapbuf_L4SB_size3 mux_bottom_track_179 (
		.in({chanx_right_in[11], bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_25_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_25_sram_inv[0:1]),
		.out(chany_bottom_out[89]));

	mux_tree_tapbuf_L4SB_size3 mux_bottom_track_181 (
		.in({chanx_right_in[9], bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_26_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_26_sram_inv[0:1]),
		.out(chany_bottom_out[90]));

	mux_tree_tapbuf_L4SB_size3 mux_bottom_track_183 (
		.in({chanx_right_in[7], bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_27_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_27_sram_inv[0:1]),
		.out(chany_bottom_out[91]));

	mux_tree_tapbuf_L4SB_size3 mux_bottom_track_185 (
		.in({chanx_right_in[5], bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_28_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_28_sram_inv[0:1]),
		.out(chany_bottom_out[92]));

	mux_tree_tapbuf_L4SB_size3 mux_bottom_track_187 (
		.in({chanx_right_in[3], bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size3_29_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_29_sram_inv[0:1]),
		.out(chany_bottom_out[93]));

	mux_tree_tapbuf_L4SB_size3_mem mem_bottom_track_63 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size4_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_0_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_0_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_bottom_track_65 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_1_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_1_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_bottom_track_77 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size4_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_2_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_2_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_bottom_track_79 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_3_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_3_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_bottom_track_91 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size4_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_4_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_4_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_bottom_track_93 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_5_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_5_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_bottom_track_105 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size4_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_6_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_6_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_bottom_track_107 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_7_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_7_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_bottom_track_119 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size4_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_8_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_8_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_bottom_track_121 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_9_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_9_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_bottom_track_137 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size2_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_10_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_10_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_bottom_track_139 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_11_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_11_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_bottom_track_141 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_12_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_12_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_bottom_track_143 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_13_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_13_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_bottom_track_145 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_14_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_14_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_bottom_track_151 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size2_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_15_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_15_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_bottom_track_153 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_16_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_16_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_bottom_track_155 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_17_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_17_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_bottom_track_157 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_18_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_18_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_bottom_track_159 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_19_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_19_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_bottom_track_165 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size2_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_20_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_20_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_bottom_track_167 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_21_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_21_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_bottom_track_169 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_22_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_22_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_bottom_track_171 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_23_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_23_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_bottom_track_173 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_24_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_24_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_bottom_track_179 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size2_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_25_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_25_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_bottom_track_181 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_26_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_26_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_bottom_track_183 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_27_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_27_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_27_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_bottom_track_185 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_27_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_28_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_28_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_28_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_bottom_track_187 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_28_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_29_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_29_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_29_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size2 mux_bottom_track_133 (
		.in({chanx_right_in[94], bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size2_0_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_0_sram_inv),
		.out(chany_bottom_out[66]));

	mux_tree_tapbuf_L4SB_size2 mux_bottom_track_135 (
		.in({chanx_right_in[90], bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size2_1_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_1_sram_inv),
		.out(chany_bottom_out[67]));

	mux_tree_tapbuf_L4SB_size2 mux_bottom_track_147 (
		.in({chanx_right_in[66], bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size2_2_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_2_sram_inv),
		.out(chany_bottom_out[73]));

	mux_tree_tapbuf_L4SB_size2 mux_bottom_track_149 (
		.in({chanx_right_in[62], bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size2_3_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_3_sram_inv),
		.out(chany_bottom_out[74]));

	mux_tree_tapbuf_L4SB_size2 mux_bottom_track_161 (
		.in({chanx_right_in[38], bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size2_4_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_4_sram_inv),
		.out(chany_bottom_out[80]));

	mux_tree_tapbuf_L4SB_size2 mux_bottom_track_163 (
		.in({chanx_right_in[34], bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size2_5_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_5_sram_inv),
		.out(chany_bottom_out[81]));

	mux_tree_tapbuf_L4SB_size2 mux_bottom_track_175 (
		.in({chanx_right_in[15], bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size2_6_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_6_sram_inv),
		.out(chany_bottom_out[87]));

	mux_tree_tapbuf_L4SB_size2 mux_bottom_track_177 (
		.in({chanx_right_in[13], bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size2_7_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_7_sram_inv),
		.out(chany_bottom_out[88]));

	mux_tree_tapbuf_L4SB_size2 mux_bottom_track_189 (
		.in({chanx_right_in[1], bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size2_8_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_8_sram_inv),
		.out(chany_bottom_out[94]));

	mux_tree_tapbuf_L4SB_size2 mux_bottom_track_191 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_, chanx_left_in[1]}),
		.sram(mux_tree_tapbuf_L4SB_size2_9_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_9_sram_inv),
		.out(chany_bottom_out[95]));

	mux_tree_tapbuf_L4SB_size2_mem mem_bottom_track_133 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size5_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size2_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size2_0_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_0_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_bottom_track_135 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size2_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size2_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size2_1_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_1_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_bottom_track_147 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size2_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size2_2_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_2_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_bottom_track_149 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size2_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size2_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size2_3_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_3_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_bottom_track_161 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size2_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size2_4_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_4_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_bottom_track_163 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size2_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size2_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size2_5_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_5_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_bottom_track_175 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size2_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size2_6_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_6_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_bottom_track_177 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size2_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size2_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size2_7_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_7_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_bottom_track_189 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_29_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size2_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size2_8_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_8_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_bottom_track_191 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size2_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size2_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size2_9_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_9_sram_inv));

	mux_tree_tapbuf_L2SB_size13 mux_left_track_5 (
		.in({chanx_right_in[2], chanx_right_in[48], chanx_right_in[88], chany_bottom_in[0], chany_bottom_in[30], chany_bottom_in[60], chany_bottom_in[90], left_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_11__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_33__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_43__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_53__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_63__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L2SB_size13_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L2SB_size13_0_sram_inv[0:3]),
		.out(chanx_left_out[2]));

	mux_tree_tapbuf_L2SB_size13 mux_left_track_9 (
		.in({chanx_right_in[4], chanx_right_in[49], chanx_right_in[89], chany_bottom_in[1], chany_bottom_in[31], chany_bottom_in[61], chany_bottom_in[91], left_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_24__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_34__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_44__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_54__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_64__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L2SB_size13_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L2SB_size13_1_sram_inv[0:3]),
		.out(chanx_left_out[4]));

	mux_tree_tapbuf_L2SB_size13 mux_left_track_13 (
		.in({chanx_right_in[6], chanx_right_in[51], chanx_right_in[91], chany_bottom_in[2], chany_bottom_in[32], chany_bottom_in[62], chany_bottom_in[92], left_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_25__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_35__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_45__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_55__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_65__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L2SB_size13_2_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L2SB_size13_2_sram_inv[0:3]),
		.out(chanx_left_out[6]));

	mux_tree_tapbuf_L2SB_size13 mux_left_track_17 (
		.in({chanx_right_in[8], chanx_right_in[52], chanx_right_in[92], chany_bottom_in[3], chany_bottom_in[33], chany_bottom_in[63], chany_bottom_in[93], left_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_26__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_36__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_46__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_56__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_66__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L2SB_size13_3_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L2SB_size13_3_sram_inv[0:3]),
		.out(chanx_left_out[8]));

	mux_tree_tapbuf_L2SB_size13 mux_left_track_21 (
		.in({chanx_right_in[10], chanx_right_in[53], chanx_right_in[93], chany_bottom_in[4], chany_bottom_in[34], chany_bottom_in[64], chany_bottom_in[94], left_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_27__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_37__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_47__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_57__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_67__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L2SB_size13_4_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L2SB_size13_4_sram_inv[0:3]),
		.out(chanx_left_out[10]));

	mux_tree_tapbuf_L2SB_size13_mem mem_left_track_5 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size12_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size13_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size13_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L2SB_size13_0_sram_inv[0:3]));

	mux_tree_tapbuf_L2SB_size13_mem mem_left_track_9 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size13_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size13_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size13_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L2SB_size13_1_sram_inv[0:3]));

	mux_tree_tapbuf_L2SB_size13_mem mem_left_track_13 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size13_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size13_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size13_2_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L2SB_size13_2_sram_inv[0:3]));

	mux_tree_tapbuf_L2SB_size13_mem mem_left_track_17 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size13_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size13_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size13_3_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L2SB_size13_3_sram_inv[0:3]));

	mux_tree_tapbuf_L2SB_size13_mem mem_left_track_21 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size13_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size13_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size13_4_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L2SB_size13_4_sram_inv[0:3]));

endmodule
// ----- END Verilog module for sb_2__8_ -----

//----- Default net type -----
`default_nettype none



