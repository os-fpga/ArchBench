//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for physical tile: io_bottom]
//	Author: Xifan TANG
//	Organization: University of Utah
//-------------------------------------------
//----- Time scale -----
`timescale 1ns / 1ps

// ----- BEGIN Grid Verilog module: grid_io_bottom -----
//----- Default net type -----
`default_nettype wire

// ----- Verilog module for grid_io_bottom -----
module grid_io_bottom(global_reset,
                      scan_mode,
                      scan_enable,
                      config_enable,
                      prog_clock,
                      gfpga_pad_RS_PREIO_A2F,
                      gfpga_pad_RS_PREIO_F2A,
                      gfpga_pad_RS_PREIO_SOC_CLK,
                      top_width_0_height_0_subtile_14__pin_f2a_i_0_,
                      top_width_0_height_0_subtile_15__pin_f2a_i_0_,
                      top_width_0_height_0_subtile_16__pin_f2a_i_0_,
                      top_width_0_height_0_subtile_17__pin_f2a_i_0_,
                      top_width_0_height_0_subtile_18__pin_f2a_i_0_,
                      top_width_0_height_0_subtile_19__pin_f2a_i_0_,
                      top_width_0_height_0_subtile_20__pin_f2a_i_0_,
                      top_width_0_height_0_subtile_21__pin_f2a_i_0_,
                      top_width_0_height_0_subtile_22__pin_f2a_i_0_,
                      top_width_0_height_0_subtile_23__pin_f2a_i_0_,
                      top_width_0_height_0_subtile_24__pin_f2a_i_0_,
                      top_width_0_height_0_subtile_25__pin_f2a_i_0_,
                      top_width_0_height_0_subtile_26__pin_f2a_i_0_,
                      top_width_0_height_0_subtile_27__pin_f2a_i_0_,
                      top_width_0_height_0_subtile_28__pin_f2a_i_0_,
                      top_width_0_height_0_subtile_29__pin_f2a_i_0_,
                      top_width_0_height_0_subtile_30__pin_f2a_i_0_,
                      top_width_0_height_0_subtile_31__pin_f2a_i_0_,
                      top_width_0_height_0_subtile_32__pin_f2a_i_0_,
                      top_width_0_height_0_subtile_33__pin_f2a_i_0_,
                      top_width_0_height_0_subtile_34__pin_f2a_i_0_,
                      top_width_0_height_0_subtile_35__pin_f2a_i_0_,
                      top_width_0_height_0_subtile_36__pin_f2a_i_0_,
                      top_width_0_height_0_subtile_37__pin_f2a_i_0_,
                      top_width_0_height_0_subtile_38__pin_f2a_i_0_,
                      top_width_0_height_0_subtile_39__pin_f2a_i_0_,
                      top_width_0_height_0_subtile_40__pin_f2a_i_0_,
                      top_width_0_height_0_subtile_41__pin_f2a_i_0_,
                      top_width_0_height_0_subtile_42__pin_f2a_i_0_,
                      top_width_0_height_0_subtile_43__pin_f2a_i_0_,
                      top_width_0_height_0_subtile_44__pin_f2a_i_0_,
                      top_width_0_height_0_subtile_45__pin_f2a_i_0_,
                      top_width_0_height_0_subtile_46__pin_f2a_i_0_,
                      top_width_0_height_0_subtile_47__pin_f2a_i_0_,
                      top_width_0_height_0_subtile_48__pin_f2a_i_0_,
                      top_width_0_height_0_subtile_49__pin_f2a_i_0_,
                      top_width_0_height_0_subtile_50__pin_f2a_i_0_,
                      top_width_0_height_0_subtile_51__pin_f2a_i_0_,
                      top_width_0_height_0_subtile_52__pin_f2a_i_0_,
                      top_width_0_height_0_subtile_53__pin_f2a_i_0_,
                      top_width_0_height_0_subtile_54__pin_f2a_i_0_,
                      top_width_0_height_0_subtile_55__pin_f2a_i_0_,
                      top_width_0_height_0_subtile_56__pin_f2a_i_0_,
                      top_width_0_height_0_subtile_57__pin_f2a_i_0_,
                      top_width_0_height_0_subtile_58__pin_f2a_i_0_,
                      top_width_0_height_0_subtile_59__pin_f2a_i_0_,
                      top_width_0_height_0_subtile_60__pin_f2a_i_0_,
                      top_width_0_height_0_subtile_61__pin_f2a_i_0_,
                      top_width_0_height_0_subtile_62__pin_f2a_i_0_,
                      top_width_0_height_0_subtile_63__pin_f2a_i_0_,
                      top_width_0_height_0_subtile_64__pin_f2a_i_0_,
                      top_width_0_height_0_subtile_65__pin_f2a_i_0_,
                      top_width_0_height_0_subtile_66__pin_f2a_i_0_,
                      top_width_0_height_0_subtile_67__pin_f2a_i_0_,
                      top_width_0_height_0_subtile_68__pin_f2a_i_0_,
                      top_width_0_height_0_subtile_69__pin_f2a_i_0_,
                      top_width_0_height_0_subtile_70__pin_f2a_i_0_,
                      top_width_0_height_0_subtile_71__pin_f2a_i_0_,
                      right_width_0_height_0_subtile_0__pin_f2a_i_0_,
                      right_width_0_height_0_subtile_1__pin_f2a_i_0_,
                      right_width_0_height_0_subtile_2__pin_f2a_i_0_,
                      right_width_0_height_0_subtile_3__pin_f2a_i_0_,
                      right_width_0_height_0_subtile_4__pin_f2a_i_0_,
                      right_width_0_height_0_subtile_5__pin_f2a_i_0_,
                      right_width_0_height_0_subtile_6__pin_f2a_i_0_,
                      right_width_0_height_0_subtile_7__pin_f2a_i_0_,
                      right_width_0_height_0_subtile_8__pin_f2a_i_0_,
                      right_width_0_height_0_subtile_9__pin_f2a_i_0_,
                      right_width_0_height_0_subtile_10__pin_f2a_i_0_,
                      right_width_0_height_0_subtile_11__pin_f2a_i_0_,
                      right_width_0_height_0_subtile_12__pin_f2a_i_0_,
                      right_width_0_height_0_subtile_13__pin_f2a_i_0_,
                      bottom_width_0_height_0_subtile_0__pin_clk_0_,
                      bottom_width_0_height_0_subtile_0__pin_clk_1_,
                      bottom_width_0_height_0_subtile_0__pin_clk_2_,
                      bottom_width_0_height_0_subtile_0__pin_clk_3_,
                      bottom_width_0_height_0_subtile_0__pin_clk_4_,
                      bottom_width_0_height_0_subtile_0__pin_clk_5_,
                      bottom_width_0_height_0_subtile_0__pin_clk_6_,
                      bottom_width_0_height_0_subtile_0__pin_clk_7_,
                      bottom_width_0_height_0_subtile_0__pin_clk_8_,
                      bottom_width_0_height_0_subtile_0__pin_clk_9_,
                      bottom_width_0_height_0_subtile_0__pin_clk_10_,
                      bottom_width_0_height_0_subtile_0__pin_clk_11_,
                      bottom_width_0_height_0_subtile_0__pin_clk_12_,
                      bottom_width_0_height_0_subtile_0__pin_clk_13_,
                      bottom_width_0_height_0_subtile_0__pin_clk_14_,
                      bottom_width_0_height_0_subtile_0__pin_clk_15_,
                      bottom_width_0_height_0_subtile_1__pin_clk_0_,
                      bottom_width_0_height_0_subtile_1__pin_clk_1_,
                      bottom_width_0_height_0_subtile_1__pin_clk_2_,
                      bottom_width_0_height_0_subtile_1__pin_clk_3_,
                      bottom_width_0_height_0_subtile_1__pin_clk_4_,
                      bottom_width_0_height_0_subtile_1__pin_clk_5_,
                      bottom_width_0_height_0_subtile_1__pin_clk_6_,
                      bottom_width_0_height_0_subtile_1__pin_clk_7_,
                      bottom_width_0_height_0_subtile_1__pin_clk_8_,
                      bottom_width_0_height_0_subtile_1__pin_clk_9_,
                      bottom_width_0_height_0_subtile_1__pin_clk_10_,
                      bottom_width_0_height_0_subtile_1__pin_clk_11_,
                      bottom_width_0_height_0_subtile_1__pin_clk_12_,
                      bottom_width_0_height_0_subtile_1__pin_clk_13_,
                      bottom_width_0_height_0_subtile_1__pin_clk_14_,
                      bottom_width_0_height_0_subtile_1__pin_clk_15_,
                      bottom_width_0_height_0_subtile_2__pin_clk_0_,
                      bottom_width_0_height_0_subtile_2__pin_clk_1_,
                      bottom_width_0_height_0_subtile_2__pin_clk_2_,
                      bottom_width_0_height_0_subtile_2__pin_clk_3_,
                      bottom_width_0_height_0_subtile_2__pin_clk_4_,
                      bottom_width_0_height_0_subtile_2__pin_clk_5_,
                      bottom_width_0_height_0_subtile_2__pin_clk_6_,
                      bottom_width_0_height_0_subtile_2__pin_clk_7_,
                      bottom_width_0_height_0_subtile_2__pin_clk_8_,
                      bottom_width_0_height_0_subtile_2__pin_clk_9_,
                      bottom_width_0_height_0_subtile_2__pin_clk_10_,
                      bottom_width_0_height_0_subtile_2__pin_clk_11_,
                      bottom_width_0_height_0_subtile_2__pin_clk_12_,
                      bottom_width_0_height_0_subtile_2__pin_clk_13_,
                      bottom_width_0_height_0_subtile_2__pin_clk_14_,
                      bottom_width_0_height_0_subtile_2__pin_clk_15_,
                      bottom_width_0_height_0_subtile_3__pin_clk_0_,
                      bottom_width_0_height_0_subtile_3__pin_clk_1_,
                      bottom_width_0_height_0_subtile_3__pin_clk_2_,
                      bottom_width_0_height_0_subtile_3__pin_clk_3_,
                      bottom_width_0_height_0_subtile_3__pin_clk_4_,
                      bottom_width_0_height_0_subtile_3__pin_clk_5_,
                      bottom_width_0_height_0_subtile_3__pin_clk_6_,
                      bottom_width_0_height_0_subtile_3__pin_clk_7_,
                      bottom_width_0_height_0_subtile_3__pin_clk_8_,
                      bottom_width_0_height_0_subtile_3__pin_clk_9_,
                      bottom_width_0_height_0_subtile_3__pin_clk_10_,
                      bottom_width_0_height_0_subtile_3__pin_clk_11_,
                      bottom_width_0_height_0_subtile_3__pin_clk_12_,
                      bottom_width_0_height_0_subtile_3__pin_clk_13_,
                      bottom_width_0_height_0_subtile_3__pin_clk_14_,
                      bottom_width_0_height_0_subtile_3__pin_clk_15_,
                      bottom_width_0_height_0_subtile_4__pin_clk_0_,
                      bottom_width_0_height_0_subtile_4__pin_clk_1_,
                      bottom_width_0_height_0_subtile_4__pin_clk_2_,
                      bottom_width_0_height_0_subtile_4__pin_clk_3_,
                      bottom_width_0_height_0_subtile_4__pin_clk_4_,
                      bottom_width_0_height_0_subtile_4__pin_clk_5_,
                      bottom_width_0_height_0_subtile_4__pin_clk_6_,
                      bottom_width_0_height_0_subtile_4__pin_clk_7_,
                      bottom_width_0_height_0_subtile_4__pin_clk_8_,
                      bottom_width_0_height_0_subtile_4__pin_clk_9_,
                      bottom_width_0_height_0_subtile_4__pin_clk_10_,
                      bottom_width_0_height_0_subtile_4__pin_clk_11_,
                      bottom_width_0_height_0_subtile_4__pin_clk_12_,
                      bottom_width_0_height_0_subtile_4__pin_clk_13_,
                      bottom_width_0_height_0_subtile_4__pin_clk_14_,
                      bottom_width_0_height_0_subtile_4__pin_clk_15_,
                      bottom_width_0_height_0_subtile_5__pin_clk_0_,
                      bottom_width_0_height_0_subtile_5__pin_clk_1_,
                      bottom_width_0_height_0_subtile_5__pin_clk_2_,
                      bottom_width_0_height_0_subtile_5__pin_clk_3_,
                      bottom_width_0_height_0_subtile_5__pin_clk_4_,
                      bottom_width_0_height_0_subtile_5__pin_clk_5_,
                      bottom_width_0_height_0_subtile_5__pin_clk_6_,
                      bottom_width_0_height_0_subtile_5__pin_clk_7_,
                      bottom_width_0_height_0_subtile_5__pin_clk_8_,
                      bottom_width_0_height_0_subtile_5__pin_clk_9_,
                      bottom_width_0_height_0_subtile_5__pin_clk_10_,
                      bottom_width_0_height_0_subtile_5__pin_clk_11_,
                      bottom_width_0_height_0_subtile_5__pin_clk_12_,
                      bottom_width_0_height_0_subtile_5__pin_clk_13_,
                      bottom_width_0_height_0_subtile_5__pin_clk_14_,
                      bottom_width_0_height_0_subtile_5__pin_clk_15_,
                      bottom_width_0_height_0_subtile_6__pin_clk_0_,
                      bottom_width_0_height_0_subtile_6__pin_clk_1_,
                      bottom_width_0_height_0_subtile_6__pin_clk_2_,
                      bottom_width_0_height_0_subtile_6__pin_clk_3_,
                      bottom_width_0_height_0_subtile_6__pin_clk_4_,
                      bottom_width_0_height_0_subtile_6__pin_clk_5_,
                      bottom_width_0_height_0_subtile_6__pin_clk_6_,
                      bottom_width_0_height_0_subtile_6__pin_clk_7_,
                      bottom_width_0_height_0_subtile_6__pin_clk_8_,
                      bottom_width_0_height_0_subtile_6__pin_clk_9_,
                      bottom_width_0_height_0_subtile_6__pin_clk_10_,
                      bottom_width_0_height_0_subtile_6__pin_clk_11_,
                      bottom_width_0_height_0_subtile_6__pin_clk_12_,
                      bottom_width_0_height_0_subtile_6__pin_clk_13_,
                      bottom_width_0_height_0_subtile_6__pin_clk_14_,
                      bottom_width_0_height_0_subtile_6__pin_clk_15_,
                      bottom_width_0_height_0_subtile_7__pin_clk_0_,
                      bottom_width_0_height_0_subtile_7__pin_clk_1_,
                      bottom_width_0_height_0_subtile_7__pin_clk_2_,
                      bottom_width_0_height_0_subtile_7__pin_clk_3_,
                      bottom_width_0_height_0_subtile_7__pin_clk_4_,
                      bottom_width_0_height_0_subtile_7__pin_clk_5_,
                      bottom_width_0_height_0_subtile_7__pin_clk_6_,
                      bottom_width_0_height_0_subtile_7__pin_clk_7_,
                      bottom_width_0_height_0_subtile_7__pin_clk_8_,
                      bottom_width_0_height_0_subtile_7__pin_clk_9_,
                      bottom_width_0_height_0_subtile_7__pin_clk_10_,
                      bottom_width_0_height_0_subtile_7__pin_clk_11_,
                      bottom_width_0_height_0_subtile_7__pin_clk_12_,
                      bottom_width_0_height_0_subtile_7__pin_clk_13_,
                      bottom_width_0_height_0_subtile_7__pin_clk_14_,
                      bottom_width_0_height_0_subtile_7__pin_clk_15_,
                      bottom_width_0_height_0_subtile_8__pin_clk_0_,
                      bottom_width_0_height_0_subtile_8__pin_clk_1_,
                      bottom_width_0_height_0_subtile_8__pin_clk_2_,
                      bottom_width_0_height_0_subtile_8__pin_clk_3_,
                      bottom_width_0_height_0_subtile_8__pin_clk_4_,
                      bottom_width_0_height_0_subtile_8__pin_clk_5_,
                      bottom_width_0_height_0_subtile_8__pin_clk_6_,
                      bottom_width_0_height_0_subtile_8__pin_clk_7_,
                      bottom_width_0_height_0_subtile_8__pin_clk_8_,
                      bottom_width_0_height_0_subtile_8__pin_clk_9_,
                      bottom_width_0_height_0_subtile_8__pin_clk_10_,
                      bottom_width_0_height_0_subtile_8__pin_clk_11_,
                      bottom_width_0_height_0_subtile_8__pin_clk_12_,
                      bottom_width_0_height_0_subtile_8__pin_clk_13_,
                      bottom_width_0_height_0_subtile_8__pin_clk_14_,
                      bottom_width_0_height_0_subtile_8__pin_clk_15_,
                      bottom_width_0_height_0_subtile_9__pin_clk_0_,
                      bottom_width_0_height_0_subtile_9__pin_clk_1_,
                      bottom_width_0_height_0_subtile_9__pin_clk_2_,
                      bottom_width_0_height_0_subtile_9__pin_clk_3_,
                      bottom_width_0_height_0_subtile_9__pin_clk_4_,
                      bottom_width_0_height_0_subtile_9__pin_clk_5_,
                      bottom_width_0_height_0_subtile_9__pin_clk_6_,
                      bottom_width_0_height_0_subtile_9__pin_clk_7_,
                      bottom_width_0_height_0_subtile_9__pin_clk_8_,
                      bottom_width_0_height_0_subtile_9__pin_clk_9_,
                      bottom_width_0_height_0_subtile_9__pin_clk_10_,
                      bottom_width_0_height_0_subtile_9__pin_clk_11_,
                      bottom_width_0_height_0_subtile_9__pin_clk_12_,
                      bottom_width_0_height_0_subtile_9__pin_clk_13_,
                      bottom_width_0_height_0_subtile_9__pin_clk_14_,
                      bottom_width_0_height_0_subtile_9__pin_clk_15_,
                      bottom_width_0_height_0_subtile_10__pin_clk_0_,
                      bottom_width_0_height_0_subtile_10__pin_clk_1_,
                      bottom_width_0_height_0_subtile_10__pin_clk_2_,
                      bottom_width_0_height_0_subtile_10__pin_clk_3_,
                      bottom_width_0_height_0_subtile_10__pin_clk_4_,
                      bottom_width_0_height_0_subtile_10__pin_clk_5_,
                      bottom_width_0_height_0_subtile_10__pin_clk_6_,
                      bottom_width_0_height_0_subtile_10__pin_clk_7_,
                      bottom_width_0_height_0_subtile_10__pin_clk_8_,
                      bottom_width_0_height_0_subtile_10__pin_clk_9_,
                      bottom_width_0_height_0_subtile_10__pin_clk_10_,
                      bottom_width_0_height_0_subtile_10__pin_clk_11_,
                      bottom_width_0_height_0_subtile_10__pin_clk_12_,
                      bottom_width_0_height_0_subtile_10__pin_clk_13_,
                      bottom_width_0_height_0_subtile_10__pin_clk_14_,
                      bottom_width_0_height_0_subtile_10__pin_clk_15_,
                      bottom_width_0_height_0_subtile_11__pin_clk_0_,
                      bottom_width_0_height_0_subtile_11__pin_clk_1_,
                      bottom_width_0_height_0_subtile_11__pin_clk_2_,
                      bottom_width_0_height_0_subtile_11__pin_clk_3_,
                      bottom_width_0_height_0_subtile_11__pin_clk_4_,
                      bottom_width_0_height_0_subtile_11__pin_clk_5_,
                      bottom_width_0_height_0_subtile_11__pin_clk_6_,
                      bottom_width_0_height_0_subtile_11__pin_clk_7_,
                      bottom_width_0_height_0_subtile_11__pin_clk_8_,
                      bottom_width_0_height_0_subtile_11__pin_clk_9_,
                      bottom_width_0_height_0_subtile_11__pin_clk_10_,
                      bottom_width_0_height_0_subtile_11__pin_clk_11_,
                      bottom_width_0_height_0_subtile_11__pin_clk_12_,
                      bottom_width_0_height_0_subtile_11__pin_clk_13_,
                      bottom_width_0_height_0_subtile_11__pin_clk_14_,
                      bottom_width_0_height_0_subtile_11__pin_clk_15_,
                      bottom_width_0_height_0_subtile_12__pin_clk_0_,
                      bottom_width_0_height_0_subtile_12__pin_clk_1_,
                      bottom_width_0_height_0_subtile_12__pin_clk_2_,
                      bottom_width_0_height_0_subtile_12__pin_clk_3_,
                      bottom_width_0_height_0_subtile_12__pin_clk_4_,
                      bottom_width_0_height_0_subtile_12__pin_clk_5_,
                      bottom_width_0_height_0_subtile_12__pin_clk_6_,
                      bottom_width_0_height_0_subtile_12__pin_clk_7_,
                      bottom_width_0_height_0_subtile_12__pin_clk_8_,
                      bottom_width_0_height_0_subtile_12__pin_clk_9_,
                      bottom_width_0_height_0_subtile_12__pin_clk_10_,
                      bottom_width_0_height_0_subtile_12__pin_clk_11_,
                      bottom_width_0_height_0_subtile_12__pin_clk_12_,
                      bottom_width_0_height_0_subtile_12__pin_clk_13_,
                      bottom_width_0_height_0_subtile_12__pin_clk_14_,
                      bottom_width_0_height_0_subtile_12__pin_clk_15_,
                      bottom_width_0_height_0_subtile_13__pin_clk_0_,
                      bottom_width_0_height_0_subtile_13__pin_clk_1_,
                      bottom_width_0_height_0_subtile_13__pin_clk_2_,
                      bottom_width_0_height_0_subtile_13__pin_clk_3_,
                      bottom_width_0_height_0_subtile_13__pin_clk_4_,
                      bottom_width_0_height_0_subtile_13__pin_clk_5_,
                      bottom_width_0_height_0_subtile_13__pin_clk_6_,
                      bottom_width_0_height_0_subtile_13__pin_clk_7_,
                      bottom_width_0_height_0_subtile_13__pin_clk_8_,
                      bottom_width_0_height_0_subtile_13__pin_clk_9_,
                      bottom_width_0_height_0_subtile_13__pin_clk_10_,
                      bottom_width_0_height_0_subtile_13__pin_clk_11_,
                      bottom_width_0_height_0_subtile_13__pin_clk_12_,
                      bottom_width_0_height_0_subtile_13__pin_clk_13_,
                      bottom_width_0_height_0_subtile_13__pin_clk_14_,
                      bottom_width_0_height_0_subtile_13__pin_clk_15_,
                      bottom_width_0_height_0_subtile_14__pin_clk_0_,
                      bottom_width_0_height_0_subtile_14__pin_clk_1_,
                      bottom_width_0_height_0_subtile_14__pin_clk_2_,
                      bottom_width_0_height_0_subtile_14__pin_clk_3_,
                      bottom_width_0_height_0_subtile_14__pin_clk_4_,
                      bottom_width_0_height_0_subtile_14__pin_clk_5_,
                      bottom_width_0_height_0_subtile_14__pin_clk_6_,
                      bottom_width_0_height_0_subtile_14__pin_clk_7_,
                      bottom_width_0_height_0_subtile_14__pin_clk_8_,
                      bottom_width_0_height_0_subtile_14__pin_clk_9_,
                      bottom_width_0_height_0_subtile_14__pin_clk_10_,
                      bottom_width_0_height_0_subtile_14__pin_clk_11_,
                      bottom_width_0_height_0_subtile_14__pin_clk_12_,
                      bottom_width_0_height_0_subtile_14__pin_clk_13_,
                      bottom_width_0_height_0_subtile_14__pin_clk_14_,
                      bottom_width_0_height_0_subtile_14__pin_clk_15_,
                      bottom_width_0_height_0_subtile_15__pin_clk_0_,
                      bottom_width_0_height_0_subtile_15__pin_clk_1_,
                      bottom_width_0_height_0_subtile_15__pin_clk_2_,
                      bottom_width_0_height_0_subtile_15__pin_clk_3_,
                      bottom_width_0_height_0_subtile_15__pin_clk_4_,
                      bottom_width_0_height_0_subtile_15__pin_clk_5_,
                      bottom_width_0_height_0_subtile_15__pin_clk_6_,
                      bottom_width_0_height_0_subtile_15__pin_clk_7_,
                      bottom_width_0_height_0_subtile_15__pin_clk_8_,
                      bottom_width_0_height_0_subtile_15__pin_clk_9_,
                      bottom_width_0_height_0_subtile_15__pin_clk_10_,
                      bottom_width_0_height_0_subtile_15__pin_clk_11_,
                      bottom_width_0_height_0_subtile_15__pin_clk_12_,
                      bottom_width_0_height_0_subtile_15__pin_clk_13_,
                      bottom_width_0_height_0_subtile_15__pin_clk_14_,
                      bottom_width_0_height_0_subtile_15__pin_clk_15_,
                      bottom_width_0_height_0_subtile_16__pin_clk_0_,
                      bottom_width_0_height_0_subtile_16__pin_clk_1_,
                      bottom_width_0_height_0_subtile_16__pin_clk_2_,
                      bottom_width_0_height_0_subtile_16__pin_clk_3_,
                      bottom_width_0_height_0_subtile_16__pin_clk_4_,
                      bottom_width_0_height_0_subtile_16__pin_clk_5_,
                      bottom_width_0_height_0_subtile_16__pin_clk_6_,
                      bottom_width_0_height_0_subtile_16__pin_clk_7_,
                      bottom_width_0_height_0_subtile_16__pin_clk_8_,
                      bottom_width_0_height_0_subtile_16__pin_clk_9_,
                      bottom_width_0_height_0_subtile_16__pin_clk_10_,
                      bottom_width_0_height_0_subtile_16__pin_clk_11_,
                      bottom_width_0_height_0_subtile_16__pin_clk_12_,
                      bottom_width_0_height_0_subtile_16__pin_clk_13_,
                      bottom_width_0_height_0_subtile_16__pin_clk_14_,
                      bottom_width_0_height_0_subtile_16__pin_clk_15_,
                      bottom_width_0_height_0_subtile_17__pin_clk_0_,
                      bottom_width_0_height_0_subtile_17__pin_clk_1_,
                      bottom_width_0_height_0_subtile_17__pin_clk_2_,
                      bottom_width_0_height_0_subtile_17__pin_clk_3_,
                      bottom_width_0_height_0_subtile_17__pin_clk_4_,
                      bottom_width_0_height_0_subtile_17__pin_clk_5_,
                      bottom_width_0_height_0_subtile_17__pin_clk_6_,
                      bottom_width_0_height_0_subtile_17__pin_clk_7_,
                      bottom_width_0_height_0_subtile_17__pin_clk_8_,
                      bottom_width_0_height_0_subtile_17__pin_clk_9_,
                      bottom_width_0_height_0_subtile_17__pin_clk_10_,
                      bottom_width_0_height_0_subtile_17__pin_clk_11_,
                      bottom_width_0_height_0_subtile_17__pin_clk_12_,
                      bottom_width_0_height_0_subtile_17__pin_clk_13_,
                      bottom_width_0_height_0_subtile_17__pin_clk_14_,
                      bottom_width_0_height_0_subtile_17__pin_clk_15_,
                      bottom_width_0_height_0_subtile_18__pin_clk_0_,
                      bottom_width_0_height_0_subtile_18__pin_clk_1_,
                      bottom_width_0_height_0_subtile_18__pin_clk_2_,
                      bottom_width_0_height_0_subtile_18__pin_clk_3_,
                      bottom_width_0_height_0_subtile_18__pin_clk_4_,
                      bottom_width_0_height_0_subtile_18__pin_clk_5_,
                      bottom_width_0_height_0_subtile_18__pin_clk_6_,
                      bottom_width_0_height_0_subtile_18__pin_clk_7_,
                      bottom_width_0_height_0_subtile_18__pin_clk_8_,
                      bottom_width_0_height_0_subtile_18__pin_clk_9_,
                      bottom_width_0_height_0_subtile_18__pin_clk_10_,
                      bottom_width_0_height_0_subtile_18__pin_clk_11_,
                      bottom_width_0_height_0_subtile_18__pin_clk_12_,
                      bottom_width_0_height_0_subtile_18__pin_clk_13_,
                      bottom_width_0_height_0_subtile_18__pin_clk_14_,
                      bottom_width_0_height_0_subtile_18__pin_clk_15_,
                      bottom_width_0_height_0_subtile_19__pin_clk_0_,
                      bottom_width_0_height_0_subtile_19__pin_clk_1_,
                      bottom_width_0_height_0_subtile_19__pin_clk_2_,
                      bottom_width_0_height_0_subtile_19__pin_clk_3_,
                      bottom_width_0_height_0_subtile_19__pin_clk_4_,
                      bottom_width_0_height_0_subtile_19__pin_clk_5_,
                      bottom_width_0_height_0_subtile_19__pin_clk_6_,
                      bottom_width_0_height_0_subtile_19__pin_clk_7_,
                      bottom_width_0_height_0_subtile_19__pin_clk_8_,
                      bottom_width_0_height_0_subtile_19__pin_clk_9_,
                      bottom_width_0_height_0_subtile_19__pin_clk_10_,
                      bottom_width_0_height_0_subtile_19__pin_clk_11_,
                      bottom_width_0_height_0_subtile_19__pin_clk_12_,
                      bottom_width_0_height_0_subtile_19__pin_clk_13_,
                      bottom_width_0_height_0_subtile_19__pin_clk_14_,
                      bottom_width_0_height_0_subtile_19__pin_clk_15_,
                      bottom_width_0_height_0_subtile_20__pin_clk_0_,
                      bottom_width_0_height_0_subtile_20__pin_clk_1_,
                      bottom_width_0_height_0_subtile_20__pin_clk_2_,
                      bottom_width_0_height_0_subtile_20__pin_clk_3_,
                      bottom_width_0_height_0_subtile_20__pin_clk_4_,
                      bottom_width_0_height_0_subtile_20__pin_clk_5_,
                      bottom_width_0_height_0_subtile_20__pin_clk_6_,
                      bottom_width_0_height_0_subtile_20__pin_clk_7_,
                      bottom_width_0_height_0_subtile_20__pin_clk_8_,
                      bottom_width_0_height_0_subtile_20__pin_clk_9_,
                      bottom_width_0_height_0_subtile_20__pin_clk_10_,
                      bottom_width_0_height_0_subtile_20__pin_clk_11_,
                      bottom_width_0_height_0_subtile_20__pin_clk_12_,
                      bottom_width_0_height_0_subtile_20__pin_clk_13_,
                      bottom_width_0_height_0_subtile_20__pin_clk_14_,
                      bottom_width_0_height_0_subtile_20__pin_clk_15_,
                      bottom_width_0_height_0_subtile_21__pin_clk_0_,
                      bottom_width_0_height_0_subtile_21__pin_clk_1_,
                      bottom_width_0_height_0_subtile_21__pin_clk_2_,
                      bottom_width_0_height_0_subtile_21__pin_clk_3_,
                      bottom_width_0_height_0_subtile_21__pin_clk_4_,
                      bottom_width_0_height_0_subtile_21__pin_clk_5_,
                      bottom_width_0_height_0_subtile_21__pin_clk_6_,
                      bottom_width_0_height_0_subtile_21__pin_clk_7_,
                      bottom_width_0_height_0_subtile_21__pin_clk_8_,
                      bottom_width_0_height_0_subtile_21__pin_clk_9_,
                      bottom_width_0_height_0_subtile_21__pin_clk_10_,
                      bottom_width_0_height_0_subtile_21__pin_clk_11_,
                      bottom_width_0_height_0_subtile_21__pin_clk_12_,
                      bottom_width_0_height_0_subtile_21__pin_clk_13_,
                      bottom_width_0_height_0_subtile_21__pin_clk_14_,
                      bottom_width_0_height_0_subtile_21__pin_clk_15_,
                      bottom_width_0_height_0_subtile_22__pin_clk_0_,
                      bottom_width_0_height_0_subtile_22__pin_clk_1_,
                      bottom_width_0_height_0_subtile_22__pin_clk_2_,
                      bottom_width_0_height_0_subtile_22__pin_clk_3_,
                      bottom_width_0_height_0_subtile_22__pin_clk_4_,
                      bottom_width_0_height_0_subtile_22__pin_clk_5_,
                      bottom_width_0_height_0_subtile_22__pin_clk_6_,
                      bottom_width_0_height_0_subtile_22__pin_clk_7_,
                      bottom_width_0_height_0_subtile_22__pin_clk_8_,
                      bottom_width_0_height_0_subtile_22__pin_clk_9_,
                      bottom_width_0_height_0_subtile_22__pin_clk_10_,
                      bottom_width_0_height_0_subtile_22__pin_clk_11_,
                      bottom_width_0_height_0_subtile_22__pin_clk_12_,
                      bottom_width_0_height_0_subtile_22__pin_clk_13_,
                      bottom_width_0_height_0_subtile_22__pin_clk_14_,
                      bottom_width_0_height_0_subtile_22__pin_clk_15_,
                      bottom_width_0_height_0_subtile_23__pin_clk_0_,
                      bottom_width_0_height_0_subtile_23__pin_clk_1_,
                      bottom_width_0_height_0_subtile_23__pin_clk_2_,
                      bottom_width_0_height_0_subtile_23__pin_clk_3_,
                      bottom_width_0_height_0_subtile_23__pin_clk_4_,
                      bottom_width_0_height_0_subtile_23__pin_clk_5_,
                      bottom_width_0_height_0_subtile_23__pin_clk_6_,
                      bottom_width_0_height_0_subtile_23__pin_clk_7_,
                      bottom_width_0_height_0_subtile_23__pin_clk_8_,
                      bottom_width_0_height_0_subtile_23__pin_clk_9_,
                      bottom_width_0_height_0_subtile_23__pin_clk_10_,
                      bottom_width_0_height_0_subtile_23__pin_clk_11_,
                      bottom_width_0_height_0_subtile_23__pin_clk_12_,
                      bottom_width_0_height_0_subtile_23__pin_clk_13_,
                      bottom_width_0_height_0_subtile_23__pin_clk_14_,
                      bottom_width_0_height_0_subtile_23__pin_clk_15_,
                      bottom_width_0_height_0_subtile_24__pin_clk_0_,
                      bottom_width_0_height_0_subtile_24__pin_clk_1_,
                      bottom_width_0_height_0_subtile_24__pin_clk_2_,
                      bottom_width_0_height_0_subtile_24__pin_clk_3_,
                      bottom_width_0_height_0_subtile_24__pin_clk_4_,
                      bottom_width_0_height_0_subtile_24__pin_clk_5_,
                      bottom_width_0_height_0_subtile_24__pin_clk_6_,
                      bottom_width_0_height_0_subtile_24__pin_clk_7_,
                      bottom_width_0_height_0_subtile_24__pin_clk_8_,
                      bottom_width_0_height_0_subtile_24__pin_clk_9_,
                      bottom_width_0_height_0_subtile_24__pin_clk_10_,
                      bottom_width_0_height_0_subtile_24__pin_clk_11_,
                      bottom_width_0_height_0_subtile_24__pin_clk_12_,
                      bottom_width_0_height_0_subtile_24__pin_clk_13_,
                      bottom_width_0_height_0_subtile_24__pin_clk_14_,
                      bottom_width_0_height_0_subtile_24__pin_clk_15_,
                      bottom_width_0_height_0_subtile_25__pin_clk_0_,
                      bottom_width_0_height_0_subtile_25__pin_clk_1_,
                      bottom_width_0_height_0_subtile_25__pin_clk_2_,
                      bottom_width_0_height_0_subtile_25__pin_clk_3_,
                      bottom_width_0_height_0_subtile_25__pin_clk_4_,
                      bottom_width_0_height_0_subtile_25__pin_clk_5_,
                      bottom_width_0_height_0_subtile_25__pin_clk_6_,
                      bottom_width_0_height_0_subtile_25__pin_clk_7_,
                      bottom_width_0_height_0_subtile_25__pin_clk_8_,
                      bottom_width_0_height_0_subtile_25__pin_clk_9_,
                      bottom_width_0_height_0_subtile_25__pin_clk_10_,
                      bottom_width_0_height_0_subtile_25__pin_clk_11_,
                      bottom_width_0_height_0_subtile_25__pin_clk_12_,
                      bottom_width_0_height_0_subtile_25__pin_clk_13_,
                      bottom_width_0_height_0_subtile_25__pin_clk_14_,
                      bottom_width_0_height_0_subtile_25__pin_clk_15_,
                      bottom_width_0_height_0_subtile_26__pin_clk_0_,
                      bottom_width_0_height_0_subtile_26__pin_clk_1_,
                      bottom_width_0_height_0_subtile_26__pin_clk_2_,
                      bottom_width_0_height_0_subtile_26__pin_clk_3_,
                      bottom_width_0_height_0_subtile_26__pin_clk_4_,
                      bottom_width_0_height_0_subtile_26__pin_clk_5_,
                      bottom_width_0_height_0_subtile_26__pin_clk_6_,
                      bottom_width_0_height_0_subtile_26__pin_clk_7_,
                      bottom_width_0_height_0_subtile_26__pin_clk_8_,
                      bottom_width_0_height_0_subtile_26__pin_clk_9_,
                      bottom_width_0_height_0_subtile_26__pin_clk_10_,
                      bottom_width_0_height_0_subtile_26__pin_clk_11_,
                      bottom_width_0_height_0_subtile_26__pin_clk_12_,
                      bottom_width_0_height_0_subtile_26__pin_clk_13_,
                      bottom_width_0_height_0_subtile_26__pin_clk_14_,
                      bottom_width_0_height_0_subtile_26__pin_clk_15_,
                      bottom_width_0_height_0_subtile_27__pin_clk_0_,
                      bottom_width_0_height_0_subtile_27__pin_clk_1_,
                      bottom_width_0_height_0_subtile_27__pin_clk_2_,
                      bottom_width_0_height_0_subtile_27__pin_clk_3_,
                      bottom_width_0_height_0_subtile_27__pin_clk_4_,
                      bottom_width_0_height_0_subtile_27__pin_clk_5_,
                      bottom_width_0_height_0_subtile_27__pin_clk_6_,
                      bottom_width_0_height_0_subtile_27__pin_clk_7_,
                      bottom_width_0_height_0_subtile_27__pin_clk_8_,
                      bottom_width_0_height_0_subtile_27__pin_clk_9_,
                      bottom_width_0_height_0_subtile_27__pin_clk_10_,
                      bottom_width_0_height_0_subtile_27__pin_clk_11_,
                      bottom_width_0_height_0_subtile_27__pin_clk_12_,
                      bottom_width_0_height_0_subtile_27__pin_clk_13_,
                      bottom_width_0_height_0_subtile_27__pin_clk_14_,
                      bottom_width_0_height_0_subtile_27__pin_clk_15_,
                      bottom_width_0_height_0_subtile_28__pin_clk_0_,
                      bottom_width_0_height_0_subtile_28__pin_clk_1_,
                      bottom_width_0_height_0_subtile_28__pin_clk_2_,
                      bottom_width_0_height_0_subtile_28__pin_clk_3_,
                      bottom_width_0_height_0_subtile_28__pin_clk_4_,
                      bottom_width_0_height_0_subtile_28__pin_clk_5_,
                      bottom_width_0_height_0_subtile_28__pin_clk_6_,
                      bottom_width_0_height_0_subtile_28__pin_clk_7_,
                      bottom_width_0_height_0_subtile_28__pin_clk_8_,
                      bottom_width_0_height_0_subtile_28__pin_clk_9_,
                      bottom_width_0_height_0_subtile_28__pin_clk_10_,
                      bottom_width_0_height_0_subtile_28__pin_clk_11_,
                      bottom_width_0_height_0_subtile_28__pin_clk_12_,
                      bottom_width_0_height_0_subtile_28__pin_clk_13_,
                      bottom_width_0_height_0_subtile_28__pin_clk_14_,
                      bottom_width_0_height_0_subtile_28__pin_clk_15_,
                      bottom_width_0_height_0_subtile_29__pin_clk_0_,
                      bottom_width_0_height_0_subtile_29__pin_clk_1_,
                      bottom_width_0_height_0_subtile_29__pin_clk_2_,
                      bottom_width_0_height_0_subtile_29__pin_clk_3_,
                      bottom_width_0_height_0_subtile_29__pin_clk_4_,
                      bottom_width_0_height_0_subtile_29__pin_clk_5_,
                      bottom_width_0_height_0_subtile_29__pin_clk_6_,
                      bottom_width_0_height_0_subtile_29__pin_clk_7_,
                      bottom_width_0_height_0_subtile_29__pin_clk_8_,
                      bottom_width_0_height_0_subtile_29__pin_clk_9_,
                      bottom_width_0_height_0_subtile_29__pin_clk_10_,
                      bottom_width_0_height_0_subtile_29__pin_clk_11_,
                      bottom_width_0_height_0_subtile_29__pin_clk_12_,
                      bottom_width_0_height_0_subtile_29__pin_clk_13_,
                      bottom_width_0_height_0_subtile_29__pin_clk_14_,
                      bottom_width_0_height_0_subtile_29__pin_clk_15_,
                      bottom_width_0_height_0_subtile_30__pin_clk_0_,
                      bottom_width_0_height_0_subtile_30__pin_clk_1_,
                      bottom_width_0_height_0_subtile_30__pin_clk_2_,
                      bottom_width_0_height_0_subtile_30__pin_clk_3_,
                      bottom_width_0_height_0_subtile_30__pin_clk_4_,
                      bottom_width_0_height_0_subtile_30__pin_clk_5_,
                      bottom_width_0_height_0_subtile_30__pin_clk_6_,
                      bottom_width_0_height_0_subtile_30__pin_clk_7_,
                      bottom_width_0_height_0_subtile_30__pin_clk_8_,
                      bottom_width_0_height_0_subtile_30__pin_clk_9_,
                      bottom_width_0_height_0_subtile_30__pin_clk_10_,
                      bottom_width_0_height_0_subtile_30__pin_clk_11_,
                      bottom_width_0_height_0_subtile_30__pin_clk_12_,
                      bottom_width_0_height_0_subtile_30__pin_clk_13_,
                      bottom_width_0_height_0_subtile_30__pin_clk_14_,
                      bottom_width_0_height_0_subtile_30__pin_clk_15_,
                      bottom_width_0_height_0_subtile_31__pin_clk_0_,
                      bottom_width_0_height_0_subtile_31__pin_clk_1_,
                      bottom_width_0_height_0_subtile_31__pin_clk_2_,
                      bottom_width_0_height_0_subtile_31__pin_clk_3_,
                      bottom_width_0_height_0_subtile_31__pin_clk_4_,
                      bottom_width_0_height_0_subtile_31__pin_clk_5_,
                      bottom_width_0_height_0_subtile_31__pin_clk_6_,
                      bottom_width_0_height_0_subtile_31__pin_clk_7_,
                      bottom_width_0_height_0_subtile_31__pin_clk_8_,
                      bottom_width_0_height_0_subtile_31__pin_clk_9_,
                      bottom_width_0_height_0_subtile_31__pin_clk_10_,
                      bottom_width_0_height_0_subtile_31__pin_clk_11_,
                      bottom_width_0_height_0_subtile_31__pin_clk_12_,
                      bottom_width_0_height_0_subtile_31__pin_clk_13_,
                      bottom_width_0_height_0_subtile_31__pin_clk_14_,
                      bottom_width_0_height_0_subtile_31__pin_clk_15_,
                      bottom_width_0_height_0_subtile_32__pin_clk_0_,
                      bottom_width_0_height_0_subtile_32__pin_clk_1_,
                      bottom_width_0_height_0_subtile_32__pin_clk_2_,
                      bottom_width_0_height_0_subtile_32__pin_clk_3_,
                      bottom_width_0_height_0_subtile_32__pin_clk_4_,
                      bottom_width_0_height_0_subtile_32__pin_clk_5_,
                      bottom_width_0_height_0_subtile_32__pin_clk_6_,
                      bottom_width_0_height_0_subtile_32__pin_clk_7_,
                      bottom_width_0_height_0_subtile_32__pin_clk_8_,
                      bottom_width_0_height_0_subtile_32__pin_clk_9_,
                      bottom_width_0_height_0_subtile_32__pin_clk_10_,
                      bottom_width_0_height_0_subtile_32__pin_clk_11_,
                      bottom_width_0_height_0_subtile_32__pin_clk_12_,
                      bottom_width_0_height_0_subtile_32__pin_clk_13_,
                      bottom_width_0_height_0_subtile_32__pin_clk_14_,
                      bottom_width_0_height_0_subtile_32__pin_clk_15_,
                      bottom_width_0_height_0_subtile_33__pin_clk_0_,
                      bottom_width_0_height_0_subtile_33__pin_clk_1_,
                      bottom_width_0_height_0_subtile_33__pin_clk_2_,
                      bottom_width_0_height_0_subtile_33__pin_clk_3_,
                      bottom_width_0_height_0_subtile_33__pin_clk_4_,
                      bottom_width_0_height_0_subtile_33__pin_clk_5_,
                      bottom_width_0_height_0_subtile_33__pin_clk_6_,
                      bottom_width_0_height_0_subtile_33__pin_clk_7_,
                      bottom_width_0_height_0_subtile_33__pin_clk_8_,
                      bottom_width_0_height_0_subtile_33__pin_clk_9_,
                      bottom_width_0_height_0_subtile_33__pin_clk_10_,
                      bottom_width_0_height_0_subtile_33__pin_clk_11_,
                      bottom_width_0_height_0_subtile_33__pin_clk_12_,
                      bottom_width_0_height_0_subtile_33__pin_clk_13_,
                      bottom_width_0_height_0_subtile_33__pin_clk_14_,
                      bottom_width_0_height_0_subtile_33__pin_clk_15_,
                      bottom_width_0_height_0_subtile_34__pin_clk_0_,
                      bottom_width_0_height_0_subtile_34__pin_clk_1_,
                      bottom_width_0_height_0_subtile_34__pin_clk_2_,
                      bottom_width_0_height_0_subtile_34__pin_clk_3_,
                      bottom_width_0_height_0_subtile_34__pin_clk_4_,
                      bottom_width_0_height_0_subtile_34__pin_clk_5_,
                      bottom_width_0_height_0_subtile_34__pin_clk_6_,
                      bottom_width_0_height_0_subtile_34__pin_clk_7_,
                      bottom_width_0_height_0_subtile_34__pin_clk_8_,
                      bottom_width_0_height_0_subtile_34__pin_clk_9_,
                      bottom_width_0_height_0_subtile_34__pin_clk_10_,
                      bottom_width_0_height_0_subtile_34__pin_clk_11_,
                      bottom_width_0_height_0_subtile_34__pin_clk_12_,
                      bottom_width_0_height_0_subtile_34__pin_clk_13_,
                      bottom_width_0_height_0_subtile_34__pin_clk_14_,
                      bottom_width_0_height_0_subtile_34__pin_clk_15_,
                      bottom_width_0_height_0_subtile_35__pin_clk_0_,
                      bottom_width_0_height_0_subtile_35__pin_clk_1_,
                      bottom_width_0_height_0_subtile_35__pin_clk_2_,
                      bottom_width_0_height_0_subtile_35__pin_clk_3_,
                      bottom_width_0_height_0_subtile_35__pin_clk_4_,
                      bottom_width_0_height_0_subtile_35__pin_clk_5_,
                      bottom_width_0_height_0_subtile_35__pin_clk_6_,
                      bottom_width_0_height_0_subtile_35__pin_clk_7_,
                      bottom_width_0_height_0_subtile_35__pin_clk_8_,
                      bottom_width_0_height_0_subtile_35__pin_clk_9_,
                      bottom_width_0_height_0_subtile_35__pin_clk_10_,
                      bottom_width_0_height_0_subtile_35__pin_clk_11_,
                      bottom_width_0_height_0_subtile_35__pin_clk_12_,
                      bottom_width_0_height_0_subtile_35__pin_clk_13_,
                      bottom_width_0_height_0_subtile_35__pin_clk_14_,
                      bottom_width_0_height_0_subtile_35__pin_clk_15_,
                      bottom_width_0_height_0_subtile_36__pin_clk_0_,
                      bottom_width_0_height_0_subtile_36__pin_clk_1_,
                      bottom_width_0_height_0_subtile_36__pin_clk_2_,
                      bottom_width_0_height_0_subtile_36__pin_clk_3_,
                      bottom_width_0_height_0_subtile_36__pin_clk_4_,
                      bottom_width_0_height_0_subtile_36__pin_clk_5_,
                      bottom_width_0_height_0_subtile_36__pin_clk_6_,
                      bottom_width_0_height_0_subtile_36__pin_clk_7_,
                      bottom_width_0_height_0_subtile_36__pin_clk_8_,
                      bottom_width_0_height_0_subtile_36__pin_clk_9_,
                      bottom_width_0_height_0_subtile_36__pin_clk_10_,
                      bottom_width_0_height_0_subtile_36__pin_clk_11_,
                      bottom_width_0_height_0_subtile_36__pin_clk_12_,
                      bottom_width_0_height_0_subtile_36__pin_clk_13_,
                      bottom_width_0_height_0_subtile_36__pin_clk_14_,
                      bottom_width_0_height_0_subtile_36__pin_clk_15_,
                      bottom_width_0_height_0_subtile_37__pin_clk_0_,
                      bottom_width_0_height_0_subtile_37__pin_clk_1_,
                      bottom_width_0_height_0_subtile_37__pin_clk_2_,
                      bottom_width_0_height_0_subtile_37__pin_clk_3_,
                      bottom_width_0_height_0_subtile_37__pin_clk_4_,
                      bottom_width_0_height_0_subtile_37__pin_clk_5_,
                      bottom_width_0_height_0_subtile_37__pin_clk_6_,
                      bottom_width_0_height_0_subtile_37__pin_clk_7_,
                      bottom_width_0_height_0_subtile_37__pin_clk_8_,
                      bottom_width_0_height_0_subtile_37__pin_clk_9_,
                      bottom_width_0_height_0_subtile_37__pin_clk_10_,
                      bottom_width_0_height_0_subtile_37__pin_clk_11_,
                      bottom_width_0_height_0_subtile_37__pin_clk_12_,
                      bottom_width_0_height_0_subtile_37__pin_clk_13_,
                      bottom_width_0_height_0_subtile_37__pin_clk_14_,
                      bottom_width_0_height_0_subtile_37__pin_clk_15_,
                      bottom_width_0_height_0_subtile_38__pin_clk_0_,
                      bottom_width_0_height_0_subtile_38__pin_clk_1_,
                      bottom_width_0_height_0_subtile_38__pin_clk_2_,
                      bottom_width_0_height_0_subtile_38__pin_clk_3_,
                      bottom_width_0_height_0_subtile_38__pin_clk_4_,
                      bottom_width_0_height_0_subtile_38__pin_clk_5_,
                      bottom_width_0_height_0_subtile_38__pin_clk_6_,
                      bottom_width_0_height_0_subtile_38__pin_clk_7_,
                      bottom_width_0_height_0_subtile_38__pin_clk_8_,
                      bottom_width_0_height_0_subtile_38__pin_clk_9_,
                      bottom_width_0_height_0_subtile_38__pin_clk_10_,
                      bottom_width_0_height_0_subtile_38__pin_clk_11_,
                      bottom_width_0_height_0_subtile_38__pin_clk_12_,
                      bottom_width_0_height_0_subtile_38__pin_clk_13_,
                      bottom_width_0_height_0_subtile_38__pin_clk_14_,
                      bottom_width_0_height_0_subtile_38__pin_clk_15_,
                      bottom_width_0_height_0_subtile_39__pin_clk_0_,
                      bottom_width_0_height_0_subtile_39__pin_clk_1_,
                      bottom_width_0_height_0_subtile_39__pin_clk_2_,
                      bottom_width_0_height_0_subtile_39__pin_clk_3_,
                      bottom_width_0_height_0_subtile_39__pin_clk_4_,
                      bottom_width_0_height_0_subtile_39__pin_clk_5_,
                      bottom_width_0_height_0_subtile_39__pin_clk_6_,
                      bottom_width_0_height_0_subtile_39__pin_clk_7_,
                      bottom_width_0_height_0_subtile_39__pin_clk_8_,
                      bottom_width_0_height_0_subtile_39__pin_clk_9_,
                      bottom_width_0_height_0_subtile_39__pin_clk_10_,
                      bottom_width_0_height_0_subtile_39__pin_clk_11_,
                      bottom_width_0_height_0_subtile_39__pin_clk_12_,
                      bottom_width_0_height_0_subtile_39__pin_clk_13_,
                      bottom_width_0_height_0_subtile_39__pin_clk_14_,
                      bottom_width_0_height_0_subtile_39__pin_clk_15_,
                      bottom_width_0_height_0_subtile_40__pin_clk_0_,
                      bottom_width_0_height_0_subtile_40__pin_clk_1_,
                      bottom_width_0_height_0_subtile_40__pin_clk_2_,
                      bottom_width_0_height_0_subtile_40__pin_clk_3_,
                      bottom_width_0_height_0_subtile_40__pin_clk_4_,
                      bottom_width_0_height_0_subtile_40__pin_clk_5_,
                      bottom_width_0_height_0_subtile_40__pin_clk_6_,
                      bottom_width_0_height_0_subtile_40__pin_clk_7_,
                      bottom_width_0_height_0_subtile_40__pin_clk_8_,
                      bottom_width_0_height_0_subtile_40__pin_clk_9_,
                      bottom_width_0_height_0_subtile_40__pin_clk_10_,
                      bottom_width_0_height_0_subtile_40__pin_clk_11_,
                      bottom_width_0_height_0_subtile_40__pin_clk_12_,
                      bottom_width_0_height_0_subtile_40__pin_clk_13_,
                      bottom_width_0_height_0_subtile_40__pin_clk_14_,
                      bottom_width_0_height_0_subtile_40__pin_clk_15_,
                      bottom_width_0_height_0_subtile_41__pin_clk_0_,
                      bottom_width_0_height_0_subtile_41__pin_clk_1_,
                      bottom_width_0_height_0_subtile_41__pin_clk_2_,
                      bottom_width_0_height_0_subtile_41__pin_clk_3_,
                      bottom_width_0_height_0_subtile_41__pin_clk_4_,
                      bottom_width_0_height_0_subtile_41__pin_clk_5_,
                      bottom_width_0_height_0_subtile_41__pin_clk_6_,
                      bottom_width_0_height_0_subtile_41__pin_clk_7_,
                      bottom_width_0_height_0_subtile_41__pin_clk_8_,
                      bottom_width_0_height_0_subtile_41__pin_clk_9_,
                      bottom_width_0_height_0_subtile_41__pin_clk_10_,
                      bottom_width_0_height_0_subtile_41__pin_clk_11_,
                      bottom_width_0_height_0_subtile_41__pin_clk_12_,
                      bottom_width_0_height_0_subtile_41__pin_clk_13_,
                      bottom_width_0_height_0_subtile_41__pin_clk_14_,
                      bottom_width_0_height_0_subtile_41__pin_clk_15_,
                      bottom_width_0_height_0_subtile_42__pin_clk_0_,
                      bottom_width_0_height_0_subtile_42__pin_clk_1_,
                      bottom_width_0_height_0_subtile_42__pin_clk_2_,
                      bottom_width_0_height_0_subtile_42__pin_clk_3_,
                      bottom_width_0_height_0_subtile_42__pin_clk_4_,
                      bottom_width_0_height_0_subtile_42__pin_clk_5_,
                      bottom_width_0_height_0_subtile_42__pin_clk_6_,
                      bottom_width_0_height_0_subtile_42__pin_clk_7_,
                      bottom_width_0_height_0_subtile_42__pin_clk_8_,
                      bottom_width_0_height_0_subtile_42__pin_clk_9_,
                      bottom_width_0_height_0_subtile_42__pin_clk_10_,
                      bottom_width_0_height_0_subtile_42__pin_clk_11_,
                      bottom_width_0_height_0_subtile_42__pin_clk_12_,
                      bottom_width_0_height_0_subtile_42__pin_clk_13_,
                      bottom_width_0_height_0_subtile_42__pin_clk_14_,
                      bottom_width_0_height_0_subtile_42__pin_clk_15_,
                      bottom_width_0_height_0_subtile_43__pin_clk_0_,
                      bottom_width_0_height_0_subtile_43__pin_clk_1_,
                      bottom_width_0_height_0_subtile_43__pin_clk_2_,
                      bottom_width_0_height_0_subtile_43__pin_clk_3_,
                      bottom_width_0_height_0_subtile_43__pin_clk_4_,
                      bottom_width_0_height_0_subtile_43__pin_clk_5_,
                      bottom_width_0_height_0_subtile_43__pin_clk_6_,
                      bottom_width_0_height_0_subtile_43__pin_clk_7_,
                      bottom_width_0_height_0_subtile_43__pin_clk_8_,
                      bottom_width_0_height_0_subtile_43__pin_clk_9_,
                      bottom_width_0_height_0_subtile_43__pin_clk_10_,
                      bottom_width_0_height_0_subtile_43__pin_clk_11_,
                      bottom_width_0_height_0_subtile_43__pin_clk_12_,
                      bottom_width_0_height_0_subtile_43__pin_clk_13_,
                      bottom_width_0_height_0_subtile_43__pin_clk_14_,
                      bottom_width_0_height_0_subtile_43__pin_clk_15_,
                      bottom_width_0_height_0_subtile_44__pin_clk_0_,
                      bottom_width_0_height_0_subtile_44__pin_clk_1_,
                      bottom_width_0_height_0_subtile_44__pin_clk_2_,
                      bottom_width_0_height_0_subtile_44__pin_clk_3_,
                      bottom_width_0_height_0_subtile_44__pin_clk_4_,
                      bottom_width_0_height_0_subtile_44__pin_clk_5_,
                      bottom_width_0_height_0_subtile_44__pin_clk_6_,
                      bottom_width_0_height_0_subtile_44__pin_clk_7_,
                      bottom_width_0_height_0_subtile_44__pin_clk_8_,
                      bottom_width_0_height_0_subtile_44__pin_clk_9_,
                      bottom_width_0_height_0_subtile_44__pin_clk_10_,
                      bottom_width_0_height_0_subtile_44__pin_clk_11_,
                      bottom_width_0_height_0_subtile_44__pin_clk_12_,
                      bottom_width_0_height_0_subtile_44__pin_clk_13_,
                      bottom_width_0_height_0_subtile_44__pin_clk_14_,
                      bottom_width_0_height_0_subtile_44__pin_clk_15_,
                      bottom_width_0_height_0_subtile_45__pin_clk_0_,
                      bottom_width_0_height_0_subtile_45__pin_clk_1_,
                      bottom_width_0_height_0_subtile_45__pin_clk_2_,
                      bottom_width_0_height_0_subtile_45__pin_clk_3_,
                      bottom_width_0_height_0_subtile_45__pin_clk_4_,
                      bottom_width_0_height_0_subtile_45__pin_clk_5_,
                      bottom_width_0_height_0_subtile_45__pin_clk_6_,
                      bottom_width_0_height_0_subtile_45__pin_clk_7_,
                      bottom_width_0_height_0_subtile_45__pin_clk_8_,
                      bottom_width_0_height_0_subtile_45__pin_clk_9_,
                      bottom_width_0_height_0_subtile_45__pin_clk_10_,
                      bottom_width_0_height_0_subtile_45__pin_clk_11_,
                      bottom_width_0_height_0_subtile_45__pin_clk_12_,
                      bottom_width_0_height_0_subtile_45__pin_clk_13_,
                      bottom_width_0_height_0_subtile_45__pin_clk_14_,
                      bottom_width_0_height_0_subtile_45__pin_clk_15_,
                      bottom_width_0_height_0_subtile_46__pin_clk_0_,
                      bottom_width_0_height_0_subtile_46__pin_clk_1_,
                      bottom_width_0_height_0_subtile_46__pin_clk_2_,
                      bottom_width_0_height_0_subtile_46__pin_clk_3_,
                      bottom_width_0_height_0_subtile_46__pin_clk_4_,
                      bottom_width_0_height_0_subtile_46__pin_clk_5_,
                      bottom_width_0_height_0_subtile_46__pin_clk_6_,
                      bottom_width_0_height_0_subtile_46__pin_clk_7_,
                      bottom_width_0_height_0_subtile_46__pin_clk_8_,
                      bottom_width_0_height_0_subtile_46__pin_clk_9_,
                      bottom_width_0_height_0_subtile_46__pin_clk_10_,
                      bottom_width_0_height_0_subtile_46__pin_clk_11_,
                      bottom_width_0_height_0_subtile_46__pin_clk_12_,
                      bottom_width_0_height_0_subtile_46__pin_clk_13_,
                      bottom_width_0_height_0_subtile_46__pin_clk_14_,
                      bottom_width_0_height_0_subtile_46__pin_clk_15_,
                      bottom_width_0_height_0_subtile_47__pin_clk_0_,
                      bottom_width_0_height_0_subtile_47__pin_clk_1_,
                      bottom_width_0_height_0_subtile_47__pin_clk_2_,
                      bottom_width_0_height_0_subtile_47__pin_clk_3_,
                      bottom_width_0_height_0_subtile_47__pin_clk_4_,
                      bottom_width_0_height_0_subtile_47__pin_clk_5_,
                      bottom_width_0_height_0_subtile_47__pin_clk_6_,
                      bottom_width_0_height_0_subtile_47__pin_clk_7_,
                      bottom_width_0_height_0_subtile_47__pin_clk_8_,
                      bottom_width_0_height_0_subtile_47__pin_clk_9_,
                      bottom_width_0_height_0_subtile_47__pin_clk_10_,
                      bottom_width_0_height_0_subtile_47__pin_clk_11_,
                      bottom_width_0_height_0_subtile_47__pin_clk_12_,
                      bottom_width_0_height_0_subtile_47__pin_clk_13_,
                      bottom_width_0_height_0_subtile_47__pin_clk_14_,
                      bottom_width_0_height_0_subtile_47__pin_clk_15_,
                      bottom_width_0_height_0_subtile_48__pin_clk_0_,
                      bottom_width_0_height_0_subtile_48__pin_clk_1_,
                      bottom_width_0_height_0_subtile_48__pin_clk_2_,
                      bottom_width_0_height_0_subtile_48__pin_clk_3_,
                      bottom_width_0_height_0_subtile_48__pin_clk_4_,
                      bottom_width_0_height_0_subtile_48__pin_clk_5_,
                      bottom_width_0_height_0_subtile_48__pin_clk_6_,
                      bottom_width_0_height_0_subtile_48__pin_clk_7_,
                      bottom_width_0_height_0_subtile_48__pin_clk_8_,
                      bottom_width_0_height_0_subtile_48__pin_clk_9_,
                      bottom_width_0_height_0_subtile_48__pin_clk_10_,
                      bottom_width_0_height_0_subtile_48__pin_clk_11_,
                      bottom_width_0_height_0_subtile_48__pin_clk_12_,
                      bottom_width_0_height_0_subtile_48__pin_clk_13_,
                      bottom_width_0_height_0_subtile_48__pin_clk_14_,
                      bottom_width_0_height_0_subtile_48__pin_clk_15_,
                      bottom_width_0_height_0_subtile_49__pin_clk_0_,
                      bottom_width_0_height_0_subtile_49__pin_clk_1_,
                      bottom_width_0_height_0_subtile_49__pin_clk_2_,
                      bottom_width_0_height_0_subtile_49__pin_clk_3_,
                      bottom_width_0_height_0_subtile_49__pin_clk_4_,
                      bottom_width_0_height_0_subtile_49__pin_clk_5_,
                      bottom_width_0_height_0_subtile_49__pin_clk_6_,
                      bottom_width_0_height_0_subtile_49__pin_clk_7_,
                      bottom_width_0_height_0_subtile_49__pin_clk_8_,
                      bottom_width_0_height_0_subtile_49__pin_clk_9_,
                      bottom_width_0_height_0_subtile_49__pin_clk_10_,
                      bottom_width_0_height_0_subtile_49__pin_clk_11_,
                      bottom_width_0_height_0_subtile_49__pin_clk_12_,
                      bottom_width_0_height_0_subtile_49__pin_clk_13_,
                      bottom_width_0_height_0_subtile_49__pin_clk_14_,
                      bottom_width_0_height_0_subtile_49__pin_clk_15_,
                      bottom_width_0_height_0_subtile_50__pin_clk_0_,
                      bottom_width_0_height_0_subtile_50__pin_clk_1_,
                      bottom_width_0_height_0_subtile_50__pin_clk_2_,
                      bottom_width_0_height_0_subtile_50__pin_clk_3_,
                      bottom_width_0_height_0_subtile_50__pin_clk_4_,
                      bottom_width_0_height_0_subtile_50__pin_clk_5_,
                      bottom_width_0_height_0_subtile_50__pin_clk_6_,
                      bottom_width_0_height_0_subtile_50__pin_clk_7_,
                      bottom_width_0_height_0_subtile_50__pin_clk_8_,
                      bottom_width_0_height_0_subtile_50__pin_clk_9_,
                      bottom_width_0_height_0_subtile_50__pin_clk_10_,
                      bottom_width_0_height_0_subtile_50__pin_clk_11_,
                      bottom_width_0_height_0_subtile_50__pin_clk_12_,
                      bottom_width_0_height_0_subtile_50__pin_clk_13_,
                      bottom_width_0_height_0_subtile_50__pin_clk_14_,
                      bottom_width_0_height_0_subtile_50__pin_clk_15_,
                      bottom_width_0_height_0_subtile_51__pin_clk_0_,
                      bottom_width_0_height_0_subtile_51__pin_clk_1_,
                      bottom_width_0_height_0_subtile_51__pin_clk_2_,
                      bottom_width_0_height_0_subtile_51__pin_clk_3_,
                      bottom_width_0_height_0_subtile_51__pin_clk_4_,
                      bottom_width_0_height_0_subtile_51__pin_clk_5_,
                      bottom_width_0_height_0_subtile_51__pin_clk_6_,
                      bottom_width_0_height_0_subtile_51__pin_clk_7_,
                      bottom_width_0_height_0_subtile_51__pin_clk_8_,
                      bottom_width_0_height_0_subtile_51__pin_clk_9_,
                      bottom_width_0_height_0_subtile_51__pin_clk_10_,
                      bottom_width_0_height_0_subtile_51__pin_clk_11_,
                      bottom_width_0_height_0_subtile_51__pin_clk_12_,
                      bottom_width_0_height_0_subtile_51__pin_clk_13_,
                      bottom_width_0_height_0_subtile_51__pin_clk_14_,
                      bottom_width_0_height_0_subtile_51__pin_clk_15_,
                      bottom_width_0_height_0_subtile_52__pin_clk_0_,
                      bottom_width_0_height_0_subtile_52__pin_clk_1_,
                      bottom_width_0_height_0_subtile_52__pin_clk_2_,
                      bottom_width_0_height_0_subtile_52__pin_clk_3_,
                      bottom_width_0_height_0_subtile_52__pin_clk_4_,
                      bottom_width_0_height_0_subtile_52__pin_clk_5_,
                      bottom_width_0_height_0_subtile_52__pin_clk_6_,
                      bottom_width_0_height_0_subtile_52__pin_clk_7_,
                      bottom_width_0_height_0_subtile_52__pin_clk_8_,
                      bottom_width_0_height_0_subtile_52__pin_clk_9_,
                      bottom_width_0_height_0_subtile_52__pin_clk_10_,
                      bottom_width_0_height_0_subtile_52__pin_clk_11_,
                      bottom_width_0_height_0_subtile_52__pin_clk_12_,
                      bottom_width_0_height_0_subtile_52__pin_clk_13_,
                      bottom_width_0_height_0_subtile_52__pin_clk_14_,
                      bottom_width_0_height_0_subtile_52__pin_clk_15_,
                      bottom_width_0_height_0_subtile_53__pin_clk_0_,
                      bottom_width_0_height_0_subtile_53__pin_clk_1_,
                      bottom_width_0_height_0_subtile_53__pin_clk_2_,
                      bottom_width_0_height_0_subtile_53__pin_clk_3_,
                      bottom_width_0_height_0_subtile_53__pin_clk_4_,
                      bottom_width_0_height_0_subtile_53__pin_clk_5_,
                      bottom_width_0_height_0_subtile_53__pin_clk_6_,
                      bottom_width_0_height_0_subtile_53__pin_clk_7_,
                      bottom_width_0_height_0_subtile_53__pin_clk_8_,
                      bottom_width_0_height_0_subtile_53__pin_clk_9_,
                      bottom_width_0_height_0_subtile_53__pin_clk_10_,
                      bottom_width_0_height_0_subtile_53__pin_clk_11_,
                      bottom_width_0_height_0_subtile_53__pin_clk_12_,
                      bottom_width_0_height_0_subtile_53__pin_clk_13_,
                      bottom_width_0_height_0_subtile_53__pin_clk_14_,
                      bottom_width_0_height_0_subtile_53__pin_clk_15_,
                      bottom_width_0_height_0_subtile_54__pin_clk_0_,
                      bottom_width_0_height_0_subtile_54__pin_clk_1_,
                      bottom_width_0_height_0_subtile_54__pin_clk_2_,
                      bottom_width_0_height_0_subtile_54__pin_clk_3_,
                      bottom_width_0_height_0_subtile_54__pin_clk_4_,
                      bottom_width_0_height_0_subtile_54__pin_clk_5_,
                      bottom_width_0_height_0_subtile_54__pin_clk_6_,
                      bottom_width_0_height_0_subtile_54__pin_clk_7_,
                      bottom_width_0_height_0_subtile_54__pin_clk_8_,
                      bottom_width_0_height_0_subtile_54__pin_clk_9_,
                      bottom_width_0_height_0_subtile_54__pin_clk_10_,
                      bottom_width_0_height_0_subtile_54__pin_clk_11_,
                      bottom_width_0_height_0_subtile_54__pin_clk_12_,
                      bottom_width_0_height_0_subtile_54__pin_clk_13_,
                      bottom_width_0_height_0_subtile_54__pin_clk_14_,
                      bottom_width_0_height_0_subtile_54__pin_clk_15_,
                      bottom_width_0_height_0_subtile_55__pin_clk_0_,
                      bottom_width_0_height_0_subtile_55__pin_clk_1_,
                      bottom_width_0_height_0_subtile_55__pin_clk_2_,
                      bottom_width_0_height_0_subtile_55__pin_clk_3_,
                      bottom_width_0_height_0_subtile_55__pin_clk_4_,
                      bottom_width_0_height_0_subtile_55__pin_clk_5_,
                      bottom_width_0_height_0_subtile_55__pin_clk_6_,
                      bottom_width_0_height_0_subtile_55__pin_clk_7_,
                      bottom_width_0_height_0_subtile_55__pin_clk_8_,
                      bottom_width_0_height_0_subtile_55__pin_clk_9_,
                      bottom_width_0_height_0_subtile_55__pin_clk_10_,
                      bottom_width_0_height_0_subtile_55__pin_clk_11_,
                      bottom_width_0_height_0_subtile_55__pin_clk_12_,
                      bottom_width_0_height_0_subtile_55__pin_clk_13_,
                      bottom_width_0_height_0_subtile_55__pin_clk_14_,
                      bottom_width_0_height_0_subtile_55__pin_clk_15_,
                      bottom_width_0_height_0_subtile_56__pin_clk_0_,
                      bottom_width_0_height_0_subtile_56__pin_clk_1_,
                      bottom_width_0_height_0_subtile_56__pin_clk_2_,
                      bottom_width_0_height_0_subtile_56__pin_clk_3_,
                      bottom_width_0_height_0_subtile_56__pin_clk_4_,
                      bottom_width_0_height_0_subtile_56__pin_clk_5_,
                      bottom_width_0_height_0_subtile_56__pin_clk_6_,
                      bottom_width_0_height_0_subtile_56__pin_clk_7_,
                      bottom_width_0_height_0_subtile_56__pin_clk_8_,
                      bottom_width_0_height_0_subtile_56__pin_clk_9_,
                      bottom_width_0_height_0_subtile_56__pin_clk_10_,
                      bottom_width_0_height_0_subtile_56__pin_clk_11_,
                      bottom_width_0_height_0_subtile_56__pin_clk_12_,
                      bottom_width_0_height_0_subtile_56__pin_clk_13_,
                      bottom_width_0_height_0_subtile_56__pin_clk_14_,
                      bottom_width_0_height_0_subtile_56__pin_clk_15_,
                      bottom_width_0_height_0_subtile_57__pin_clk_0_,
                      bottom_width_0_height_0_subtile_57__pin_clk_1_,
                      bottom_width_0_height_0_subtile_57__pin_clk_2_,
                      bottom_width_0_height_0_subtile_57__pin_clk_3_,
                      bottom_width_0_height_0_subtile_57__pin_clk_4_,
                      bottom_width_0_height_0_subtile_57__pin_clk_5_,
                      bottom_width_0_height_0_subtile_57__pin_clk_6_,
                      bottom_width_0_height_0_subtile_57__pin_clk_7_,
                      bottom_width_0_height_0_subtile_57__pin_clk_8_,
                      bottom_width_0_height_0_subtile_57__pin_clk_9_,
                      bottom_width_0_height_0_subtile_57__pin_clk_10_,
                      bottom_width_0_height_0_subtile_57__pin_clk_11_,
                      bottom_width_0_height_0_subtile_57__pin_clk_12_,
                      bottom_width_0_height_0_subtile_57__pin_clk_13_,
                      bottom_width_0_height_0_subtile_57__pin_clk_14_,
                      bottom_width_0_height_0_subtile_57__pin_clk_15_,
                      bottom_width_0_height_0_subtile_58__pin_clk_0_,
                      bottom_width_0_height_0_subtile_58__pin_clk_1_,
                      bottom_width_0_height_0_subtile_58__pin_clk_2_,
                      bottom_width_0_height_0_subtile_58__pin_clk_3_,
                      bottom_width_0_height_0_subtile_58__pin_clk_4_,
                      bottom_width_0_height_0_subtile_58__pin_clk_5_,
                      bottom_width_0_height_0_subtile_58__pin_clk_6_,
                      bottom_width_0_height_0_subtile_58__pin_clk_7_,
                      bottom_width_0_height_0_subtile_58__pin_clk_8_,
                      bottom_width_0_height_0_subtile_58__pin_clk_9_,
                      bottom_width_0_height_0_subtile_58__pin_clk_10_,
                      bottom_width_0_height_0_subtile_58__pin_clk_11_,
                      bottom_width_0_height_0_subtile_58__pin_clk_12_,
                      bottom_width_0_height_0_subtile_58__pin_clk_13_,
                      bottom_width_0_height_0_subtile_58__pin_clk_14_,
                      bottom_width_0_height_0_subtile_58__pin_clk_15_,
                      bottom_width_0_height_0_subtile_59__pin_clk_0_,
                      bottom_width_0_height_0_subtile_59__pin_clk_1_,
                      bottom_width_0_height_0_subtile_59__pin_clk_2_,
                      bottom_width_0_height_0_subtile_59__pin_clk_3_,
                      bottom_width_0_height_0_subtile_59__pin_clk_4_,
                      bottom_width_0_height_0_subtile_59__pin_clk_5_,
                      bottom_width_0_height_0_subtile_59__pin_clk_6_,
                      bottom_width_0_height_0_subtile_59__pin_clk_7_,
                      bottom_width_0_height_0_subtile_59__pin_clk_8_,
                      bottom_width_0_height_0_subtile_59__pin_clk_9_,
                      bottom_width_0_height_0_subtile_59__pin_clk_10_,
                      bottom_width_0_height_0_subtile_59__pin_clk_11_,
                      bottom_width_0_height_0_subtile_59__pin_clk_12_,
                      bottom_width_0_height_0_subtile_59__pin_clk_13_,
                      bottom_width_0_height_0_subtile_59__pin_clk_14_,
                      bottom_width_0_height_0_subtile_59__pin_clk_15_,
                      bottom_width_0_height_0_subtile_60__pin_clk_0_,
                      bottom_width_0_height_0_subtile_60__pin_clk_1_,
                      bottom_width_0_height_0_subtile_60__pin_clk_2_,
                      bottom_width_0_height_0_subtile_60__pin_clk_3_,
                      bottom_width_0_height_0_subtile_60__pin_clk_4_,
                      bottom_width_0_height_0_subtile_60__pin_clk_5_,
                      bottom_width_0_height_0_subtile_60__pin_clk_6_,
                      bottom_width_0_height_0_subtile_60__pin_clk_7_,
                      bottom_width_0_height_0_subtile_60__pin_clk_8_,
                      bottom_width_0_height_0_subtile_60__pin_clk_9_,
                      bottom_width_0_height_0_subtile_60__pin_clk_10_,
                      bottom_width_0_height_0_subtile_60__pin_clk_11_,
                      bottom_width_0_height_0_subtile_60__pin_clk_12_,
                      bottom_width_0_height_0_subtile_60__pin_clk_13_,
                      bottom_width_0_height_0_subtile_60__pin_clk_14_,
                      bottom_width_0_height_0_subtile_60__pin_clk_15_,
                      bottom_width_0_height_0_subtile_61__pin_clk_0_,
                      bottom_width_0_height_0_subtile_61__pin_clk_1_,
                      bottom_width_0_height_0_subtile_61__pin_clk_2_,
                      bottom_width_0_height_0_subtile_61__pin_clk_3_,
                      bottom_width_0_height_0_subtile_61__pin_clk_4_,
                      bottom_width_0_height_0_subtile_61__pin_clk_5_,
                      bottom_width_0_height_0_subtile_61__pin_clk_6_,
                      bottom_width_0_height_0_subtile_61__pin_clk_7_,
                      bottom_width_0_height_0_subtile_61__pin_clk_8_,
                      bottom_width_0_height_0_subtile_61__pin_clk_9_,
                      bottom_width_0_height_0_subtile_61__pin_clk_10_,
                      bottom_width_0_height_0_subtile_61__pin_clk_11_,
                      bottom_width_0_height_0_subtile_61__pin_clk_12_,
                      bottom_width_0_height_0_subtile_61__pin_clk_13_,
                      bottom_width_0_height_0_subtile_61__pin_clk_14_,
                      bottom_width_0_height_0_subtile_61__pin_clk_15_,
                      bottom_width_0_height_0_subtile_62__pin_clk_0_,
                      bottom_width_0_height_0_subtile_62__pin_clk_1_,
                      bottom_width_0_height_0_subtile_62__pin_clk_2_,
                      bottom_width_0_height_0_subtile_62__pin_clk_3_,
                      bottom_width_0_height_0_subtile_62__pin_clk_4_,
                      bottom_width_0_height_0_subtile_62__pin_clk_5_,
                      bottom_width_0_height_0_subtile_62__pin_clk_6_,
                      bottom_width_0_height_0_subtile_62__pin_clk_7_,
                      bottom_width_0_height_0_subtile_62__pin_clk_8_,
                      bottom_width_0_height_0_subtile_62__pin_clk_9_,
                      bottom_width_0_height_0_subtile_62__pin_clk_10_,
                      bottom_width_0_height_0_subtile_62__pin_clk_11_,
                      bottom_width_0_height_0_subtile_62__pin_clk_12_,
                      bottom_width_0_height_0_subtile_62__pin_clk_13_,
                      bottom_width_0_height_0_subtile_62__pin_clk_14_,
                      bottom_width_0_height_0_subtile_62__pin_clk_15_,
                      bottom_width_0_height_0_subtile_63__pin_clk_0_,
                      bottom_width_0_height_0_subtile_63__pin_clk_1_,
                      bottom_width_0_height_0_subtile_63__pin_clk_2_,
                      bottom_width_0_height_0_subtile_63__pin_clk_3_,
                      bottom_width_0_height_0_subtile_63__pin_clk_4_,
                      bottom_width_0_height_0_subtile_63__pin_clk_5_,
                      bottom_width_0_height_0_subtile_63__pin_clk_6_,
                      bottom_width_0_height_0_subtile_63__pin_clk_7_,
                      bottom_width_0_height_0_subtile_63__pin_clk_8_,
                      bottom_width_0_height_0_subtile_63__pin_clk_9_,
                      bottom_width_0_height_0_subtile_63__pin_clk_10_,
                      bottom_width_0_height_0_subtile_63__pin_clk_11_,
                      bottom_width_0_height_0_subtile_63__pin_clk_12_,
                      bottom_width_0_height_0_subtile_63__pin_clk_13_,
                      bottom_width_0_height_0_subtile_63__pin_clk_14_,
                      bottom_width_0_height_0_subtile_63__pin_clk_15_,
                      bottom_width_0_height_0_subtile_64__pin_clk_0_,
                      bottom_width_0_height_0_subtile_64__pin_clk_1_,
                      bottom_width_0_height_0_subtile_64__pin_clk_2_,
                      bottom_width_0_height_0_subtile_64__pin_clk_3_,
                      bottom_width_0_height_0_subtile_64__pin_clk_4_,
                      bottom_width_0_height_0_subtile_64__pin_clk_5_,
                      bottom_width_0_height_0_subtile_64__pin_clk_6_,
                      bottom_width_0_height_0_subtile_64__pin_clk_7_,
                      bottom_width_0_height_0_subtile_64__pin_clk_8_,
                      bottom_width_0_height_0_subtile_64__pin_clk_9_,
                      bottom_width_0_height_0_subtile_64__pin_clk_10_,
                      bottom_width_0_height_0_subtile_64__pin_clk_11_,
                      bottom_width_0_height_0_subtile_64__pin_clk_12_,
                      bottom_width_0_height_0_subtile_64__pin_clk_13_,
                      bottom_width_0_height_0_subtile_64__pin_clk_14_,
                      bottom_width_0_height_0_subtile_64__pin_clk_15_,
                      bottom_width_0_height_0_subtile_65__pin_clk_0_,
                      bottom_width_0_height_0_subtile_65__pin_clk_1_,
                      bottom_width_0_height_0_subtile_65__pin_clk_2_,
                      bottom_width_0_height_0_subtile_65__pin_clk_3_,
                      bottom_width_0_height_0_subtile_65__pin_clk_4_,
                      bottom_width_0_height_0_subtile_65__pin_clk_5_,
                      bottom_width_0_height_0_subtile_65__pin_clk_6_,
                      bottom_width_0_height_0_subtile_65__pin_clk_7_,
                      bottom_width_0_height_0_subtile_65__pin_clk_8_,
                      bottom_width_0_height_0_subtile_65__pin_clk_9_,
                      bottom_width_0_height_0_subtile_65__pin_clk_10_,
                      bottom_width_0_height_0_subtile_65__pin_clk_11_,
                      bottom_width_0_height_0_subtile_65__pin_clk_12_,
                      bottom_width_0_height_0_subtile_65__pin_clk_13_,
                      bottom_width_0_height_0_subtile_65__pin_clk_14_,
                      bottom_width_0_height_0_subtile_65__pin_clk_15_,
                      bottom_width_0_height_0_subtile_66__pin_clk_0_,
                      bottom_width_0_height_0_subtile_66__pin_clk_1_,
                      bottom_width_0_height_0_subtile_66__pin_clk_2_,
                      bottom_width_0_height_0_subtile_66__pin_clk_3_,
                      bottom_width_0_height_0_subtile_66__pin_clk_4_,
                      bottom_width_0_height_0_subtile_66__pin_clk_5_,
                      bottom_width_0_height_0_subtile_66__pin_clk_6_,
                      bottom_width_0_height_0_subtile_66__pin_clk_7_,
                      bottom_width_0_height_0_subtile_66__pin_clk_8_,
                      bottom_width_0_height_0_subtile_66__pin_clk_9_,
                      bottom_width_0_height_0_subtile_66__pin_clk_10_,
                      bottom_width_0_height_0_subtile_66__pin_clk_11_,
                      bottom_width_0_height_0_subtile_66__pin_clk_12_,
                      bottom_width_0_height_0_subtile_66__pin_clk_13_,
                      bottom_width_0_height_0_subtile_66__pin_clk_14_,
                      bottom_width_0_height_0_subtile_66__pin_clk_15_,
                      bottom_width_0_height_0_subtile_67__pin_clk_0_,
                      bottom_width_0_height_0_subtile_67__pin_clk_1_,
                      bottom_width_0_height_0_subtile_67__pin_clk_2_,
                      bottom_width_0_height_0_subtile_67__pin_clk_3_,
                      bottom_width_0_height_0_subtile_67__pin_clk_4_,
                      bottom_width_0_height_0_subtile_67__pin_clk_5_,
                      bottom_width_0_height_0_subtile_67__pin_clk_6_,
                      bottom_width_0_height_0_subtile_67__pin_clk_7_,
                      bottom_width_0_height_0_subtile_67__pin_clk_8_,
                      bottom_width_0_height_0_subtile_67__pin_clk_9_,
                      bottom_width_0_height_0_subtile_67__pin_clk_10_,
                      bottom_width_0_height_0_subtile_67__pin_clk_11_,
                      bottom_width_0_height_0_subtile_67__pin_clk_12_,
                      bottom_width_0_height_0_subtile_67__pin_clk_13_,
                      bottom_width_0_height_0_subtile_67__pin_clk_14_,
                      bottom_width_0_height_0_subtile_67__pin_clk_15_,
                      bottom_width_0_height_0_subtile_68__pin_clk_0_,
                      bottom_width_0_height_0_subtile_68__pin_clk_1_,
                      bottom_width_0_height_0_subtile_68__pin_clk_2_,
                      bottom_width_0_height_0_subtile_68__pin_clk_3_,
                      bottom_width_0_height_0_subtile_68__pin_clk_4_,
                      bottom_width_0_height_0_subtile_68__pin_clk_5_,
                      bottom_width_0_height_0_subtile_68__pin_clk_6_,
                      bottom_width_0_height_0_subtile_68__pin_clk_7_,
                      bottom_width_0_height_0_subtile_68__pin_clk_8_,
                      bottom_width_0_height_0_subtile_68__pin_clk_9_,
                      bottom_width_0_height_0_subtile_68__pin_clk_10_,
                      bottom_width_0_height_0_subtile_68__pin_clk_11_,
                      bottom_width_0_height_0_subtile_68__pin_clk_12_,
                      bottom_width_0_height_0_subtile_68__pin_clk_13_,
                      bottom_width_0_height_0_subtile_68__pin_clk_14_,
                      bottom_width_0_height_0_subtile_68__pin_clk_15_,
                      bottom_width_0_height_0_subtile_69__pin_clk_0_,
                      bottom_width_0_height_0_subtile_69__pin_clk_1_,
                      bottom_width_0_height_0_subtile_69__pin_clk_2_,
                      bottom_width_0_height_0_subtile_69__pin_clk_3_,
                      bottom_width_0_height_0_subtile_69__pin_clk_4_,
                      bottom_width_0_height_0_subtile_69__pin_clk_5_,
                      bottom_width_0_height_0_subtile_69__pin_clk_6_,
                      bottom_width_0_height_0_subtile_69__pin_clk_7_,
                      bottom_width_0_height_0_subtile_69__pin_clk_8_,
                      bottom_width_0_height_0_subtile_69__pin_clk_9_,
                      bottom_width_0_height_0_subtile_69__pin_clk_10_,
                      bottom_width_0_height_0_subtile_69__pin_clk_11_,
                      bottom_width_0_height_0_subtile_69__pin_clk_12_,
                      bottom_width_0_height_0_subtile_69__pin_clk_13_,
                      bottom_width_0_height_0_subtile_69__pin_clk_14_,
                      bottom_width_0_height_0_subtile_69__pin_clk_15_,
                      bottom_width_0_height_0_subtile_70__pin_clk_0_,
                      bottom_width_0_height_0_subtile_70__pin_clk_1_,
                      bottom_width_0_height_0_subtile_70__pin_clk_2_,
                      bottom_width_0_height_0_subtile_70__pin_clk_3_,
                      bottom_width_0_height_0_subtile_70__pin_clk_4_,
                      bottom_width_0_height_0_subtile_70__pin_clk_5_,
                      bottom_width_0_height_0_subtile_70__pin_clk_6_,
                      bottom_width_0_height_0_subtile_70__pin_clk_7_,
                      bottom_width_0_height_0_subtile_70__pin_clk_8_,
                      bottom_width_0_height_0_subtile_70__pin_clk_9_,
                      bottom_width_0_height_0_subtile_70__pin_clk_10_,
                      bottom_width_0_height_0_subtile_70__pin_clk_11_,
                      bottom_width_0_height_0_subtile_70__pin_clk_12_,
                      bottom_width_0_height_0_subtile_70__pin_clk_13_,
                      bottom_width_0_height_0_subtile_70__pin_clk_14_,
                      bottom_width_0_height_0_subtile_70__pin_clk_15_,
                      bottom_width_0_height_0_subtile_71__pin_clk_0_,
                      bottom_width_0_height_0_subtile_71__pin_clk_1_,
                      bottom_width_0_height_0_subtile_71__pin_clk_2_,
                      bottom_width_0_height_0_subtile_71__pin_clk_3_,
                      bottom_width_0_height_0_subtile_71__pin_clk_4_,
                      bottom_width_0_height_0_subtile_71__pin_clk_5_,
                      bottom_width_0_height_0_subtile_71__pin_clk_6_,
                      bottom_width_0_height_0_subtile_71__pin_clk_7_,
                      bottom_width_0_height_0_subtile_71__pin_clk_8_,
                      bottom_width_0_height_0_subtile_71__pin_clk_9_,
                      bottom_width_0_height_0_subtile_71__pin_clk_10_,
                      bottom_width_0_height_0_subtile_71__pin_clk_11_,
                      bottom_width_0_height_0_subtile_71__pin_clk_12_,
                      bottom_width_0_height_0_subtile_71__pin_clk_13_,
                      bottom_width_0_height_0_subtile_71__pin_clk_14_,
                      bottom_width_0_height_0_subtile_71__pin_clk_15_,
                      left_width_0_height_0_subtile_0__pin_sc_in_0_,
                      left_width_0_height_0_subtile_1__pin_sc_in_0_,
                      left_width_0_height_0_subtile_2__pin_sc_in_0_,
                      left_width_0_height_0_subtile_3__pin_sc_in_0_,
                      left_width_0_height_0_subtile_4__pin_sc_in_0_,
                      left_width_0_height_0_subtile_5__pin_sc_in_0_,
                      left_width_0_height_0_subtile_6__pin_sc_in_0_,
                      left_width_0_height_0_subtile_7__pin_sc_in_0_,
                      left_width_0_height_0_subtile_8__pin_sc_in_0_,
                      left_width_0_height_0_subtile_9__pin_sc_in_0_,
                      left_width_0_height_0_subtile_10__pin_sc_in_0_,
                      left_width_0_height_0_subtile_11__pin_sc_in_0_,
                      left_width_0_height_0_subtile_12__pin_sc_in_0_,
                      left_width_0_height_0_subtile_13__pin_sc_in_0_,
                      left_width_0_height_0_subtile_14__pin_sc_in_0_,
                      left_width_0_height_0_subtile_15__pin_sc_in_0_,
                      left_width_0_height_0_subtile_16__pin_sc_in_0_,
                      left_width_0_height_0_subtile_17__pin_sc_in_0_,
                      left_width_0_height_0_subtile_18__pin_sc_in_0_,
                      left_width_0_height_0_subtile_19__pin_sc_in_0_,
                      left_width_0_height_0_subtile_20__pin_sc_in_0_,
                      left_width_0_height_0_subtile_21__pin_sc_in_0_,
                      left_width_0_height_0_subtile_22__pin_sc_in_0_,
                      left_width_0_height_0_subtile_23__pin_sc_in_0_,
                      left_width_0_height_0_subtile_24__pin_sc_in_0_,
                      left_width_0_height_0_subtile_25__pin_sc_in_0_,
                      left_width_0_height_0_subtile_26__pin_sc_in_0_,
                      left_width_0_height_0_subtile_27__pin_sc_in_0_,
                      left_width_0_height_0_subtile_28__pin_sc_in_0_,
                      left_width_0_height_0_subtile_29__pin_sc_in_0_,
                      left_width_0_height_0_subtile_30__pin_sc_in_0_,
                      left_width_0_height_0_subtile_31__pin_sc_in_0_,
                      left_width_0_height_0_subtile_32__pin_sc_in_0_,
                      left_width_0_height_0_subtile_33__pin_sc_in_0_,
                      left_width_0_height_0_subtile_34__pin_sc_in_0_,
                      left_width_0_height_0_subtile_35__pin_sc_in_0_,
                      left_width_0_height_0_subtile_36__pin_sc_in_0_,
                      left_width_0_height_0_subtile_37__pin_sc_in_0_,
                      left_width_0_height_0_subtile_38__pin_sc_in_0_,
                      left_width_0_height_0_subtile_39__pin_sc_in_0_,
                      left_width_0_height_0_subtile_40__pin_sc_in_0_,
                      left_width_0_height_0_subtile_41__pin_sc_in_0_,
                      left_width_0_height_0_subtile_42__pin_sc_in_0_,
                      left_width_0_height_0_subtile_43__pin_sc_in_0_,
                      left_width_0_height_0_subtile_44__pin_sc_in_0_,
                      left_width_0_height_0_subtile_45__pin_sc_in_0_,
                      left_width_0_height_0_subtile_46__pin_sc_in_0_,
                      left_width_0_height_0_subtile_47__pin_sc_in_0_,
                      left_width_0_height_0_subtile_48__pin_sc_in_0_,
                      left_width_0_height_0_subtile_49__pin_sc_in_0_,
                      left_width_0_height_0_subtile_50__pin_sc_in_0_,
                      left_width_0_height_0_subtile_51__pin_sc_in_0_,
                      left_width_0_height_0_subtile_52__pin_sc_in_0_,
                      left_width_0_height_0_subtile_53__pin_sc_in_0_,
                      left_width_0_height_0_subtile_54__pin_sc_in_0_,
                      left_width_0_height_0_subtile_55__pin_sc_in_0_,
                      left_width_0_height_0_subtile_56__pin_sc_in_0_,
                      left_width_0_height_0_subtile_57__pin_sc_in_0_,
                      left_width_0_height_0_subtile_58__pin_sc_in_0_,
                      left_width_0_height_0_subtile_59__pin_sc_in_0_,
                      left_width_0_height_0_subtile_60__pin_sc_in_0_,
                      left_width_0_height_0_subtile_61__pin_sc_in_0_,
                      left_width_0_height_0_subtile_62__pin_sc_in_0_,
                      left_width_0_height_0_subtile_63__pin_sc_in_0_,
                      left_width_0_height_0_subtile_64__pin_sc_in_0_,
                      left_width_0_height_0_subtile_65__pin_sc_in_0_,
                      left_width_0_height_0_subtile_66__pin_sc_in_0_,
                      left_width_0_height_0_subtile_67__pin_sc_in_0_,
                      left_width_0_height_0_subtile_68__pin_sc_in_0_,
                      left_width_0_height_0_subtile_69__pin_sc_in_0_,
                      left_width_0_height_0_subtile_70__pin_sc_in_0_,
                      left_width_0_height_0_subtile_71__pin_sc_in_0_,
                      ccff_head,
                      right_width_0_height_0_subtile_12__pin_a2f_o_0_,
                      right_width_0_height_0_subtile_13__pin_a2f_o_0_,
                      right_width_0_height_0_subtile_14__pin_a2f_o_0_,
                      right_width_0_height_0_subtile_15__pin_a2f_o_0_,
                      right_width_0_height_0_subtile_16__pin_a2f_o_0_,
                      right_width_0_height_0_subtile_17__pin_a2f_o_0_,
                      right_width_0_height_0_subtile_18__pin_a2f_o_0_,
                      right_width_0_height_0_subtile_19__pin_a2f_o_0_,
                      right_width_0_height_0_subtile_20__pin_a2f_o_0_,
                      right_width_0_height_0_subtile_21__pin_a2f_o_0_,
                      right_width_0_height_0_subtile_22__pin_a2f_o_0_,
                      right_width_0_height_0_subtile_23__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_0__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_1__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_2__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_3__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_4__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_5__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_6__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_7__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_8__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_9__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_10__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_11__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_24__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_25__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_26__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_27__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_28__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_29__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_30__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_31__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_32__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_33__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_34__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_35__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_36__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_37__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_38__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_39__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_40__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_41__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_42__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_43__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_44__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_45__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_46__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_47__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_48__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_49__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_50__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_51__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_52__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_53__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_54__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_55__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_56__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_57__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_58__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_59__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_60__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_61__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_62__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_63__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_64__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_65__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_66__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_67__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_68__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_69__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_70__pin_a2f_o_0_,
                      bottom_width_0_height_0_subtile_71__pin_a2f_o_0_,
                      left_width_0_height_0_subtile_0__pin_sc_out_0_,
                      left_width_0_height_0_subtile_1__pin_sc_out_0_,
                      left_width_0_height_0_subtile_2__pin_sc_out_0_,
                      left_width_0_height_0_subtile_3__pin_sc_out_0_,
                      left_width_0_height_0_subtile_4__pin_sc_out_0_,
                      left_width_0_height_0_subtile_5__pin_sc_out_0_,
                      left_width_0_height_0_subtile_6__pin_sc_out_0_,
                      left_width_0_height_0_subtile_7__pin_sc_out_0_,
                      left_width_0_height_0_subtile_8__pin_sc_out_0_,
                      left_width_0_height_0_subtile_9__pin_sc_out_0_,
                      left_width_0_height_0_subtile_10__pin_sc_out_0_,
                      left_width_0_height_0_subtile_11__pin_sc_out_0_,
                      left_width_0_height_0_subtile_12__pin_sc_out_0_,
                      left_width_0_height_0_subtile_13__pin_sc_out_0_,
                      left_width_0_height_0_subtile_14__pin_sc_out_0_,
                      left_width_0_height_0_subtile_15__pin_sc_out_0_,
                      left_width_0_height_0_subtile_16__pin_sc_out_0_,
                      left_width_0_height_0_subtile_17__pin_sc_out_0_,
                      left_width_0_height_0_subtile_18__pin_sc_out_0_,
                      left_width_0_height_0_subtile_19__pin_sc_out_0_,
                      left_width_0_height_0_subtile_20__pin_sc_out_0_,
                      left_width_0_height_0_subtile_21__pin_sc_out_0_,
                      left_width_0_height_0_subtile_22__pin_sc_out_0_,
                      left_width_0_height_0_subtile_23__pin_sc_out_0_,
                      left_width_0_height_0_subtile_24__pin_sc_out_0_,
                      left_width_0_height_0_subtile_25__pin_sc_out_0_,
                      left_width_0_height_0_subtile_26__pin_sc_out_0_,
                      left_width_0_height_0_subtile_27__pin_sc_out_0_,
                      left_width_0_height_0_subtile_28__pin_sc_out_0_,
                      left_width_0_height_0_subtile_29__pin_sc_out_0_,
                      left_width_0_height_0_subtile_30__pin_sc_out_0_,
                      left_width_0_height_0_subtile_31__pin_sc_out_0_,
                      left_width_0_height_0_subtile_32__pin_sc_out_0_,
                      left_width_0_height_0_subtile_33__pin_sc_out_0_,
                      left_width_0_height_0_subtile_34__pin_sc_out_0_,
                      left_width_0_height_0_subtile_35__pin_sc_out_0_,
                      left_width_0_height_0_subtile_36__pin_sc_out_0_,
                      left_width_0_height_0_subtile_37__pin_sc_out_0_,
                      left_width_0_height_0_subtile_38__pin_sc_out_0_,
                      left_width_0_height_0_subtile_39__pin_sc_out_0_,
                      left_width_0_height_0_subtile_40__pin_sc_out_0_,
                      left_width_0_height_0_subtile_41__pin_sc_out_0_,
                      left_width_0_height_0_subtile_42__pin_sc_out_0_,
                      left_width_0_height_0_subtile_43__pin_sc_out_0_,
                      left_width_0_height_0_subtile_44__pin_sc_out_0_,
                      left_width_0_height_0_subtile_45__pin_sc_out_0_,
                      left_width_0_height_0_subtile_46__pin_sc_out_0_,
                      left_width_0_height_0_subtile_47__pin_sc_out_0_,
                      left_width_0_height_0_subtile_48__pin_sc_out_0_,
                      left_width_0_height_0_subtile_49__pin_sc_out_0_,
                      left_width_0_height_0_subtile_50__pin_sc_out_0_,
                      left_width_0_height_0_subtile_51__pin_sc_out_0_,
                      left_width_0_height_0_subtile_52__pin_sc_out_0_,
                      left_width_0_height_0_subtile_53__pin_sc_out_0_,
                      left_width_0_height_0_subtile_54__pin_sc_out_0_,
                      left_width_0_height_0_subtile_55__pin_sc_out_0_,
                      left_width_0_height_0_subtile_56__pin_sc_out_0_,
                      left_width_0_height_0_subtile_57__pin_sc_out_0_,
                      left_width_0_height_0_subtile_58__pin_sc_out_0_,
                      left_width_0_height_0_subtile_59__pin_sc_out_0_,
                      left_width_0_height_0_subtile_60__pin_sc_out_0_,
                      left_width_0_height_0_subtile_61__pin_sc_out_0_,
                      left_width_0_height_0_subtile_62__pin_sc_out_0_,
                      left_width_0_height_0_subtile_63__pin_sc_out_0_,
                      left_width_0_height_0_subtile_64__pin_sc_out_0_,
                      left_width_0_height_0_subtile_65__pin_sc_out_0_,
                      left_width_0_height_0_subtile_66__pin_sc_out_0_,
                      left_width_0_height_0_subtile_67__pin_sc_out_0_,
                      left_width_0_height_0_subtile_68__pin_sc_out_0_,
                      left_width_0_height_0_subtile_69__pin_sc_out_0_,
                      left_width_0_height_0_subtile_70__pin_sc_out_0_,
                      left_width_0_height_0_subtile_71__pin_sc_out_0_,
                      ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] global_reset;
//----- GLOBAL PORTS -----
input [0:0] scan_mode;
//----- GLOBAL PORTS -----
input [0:0] scan_enable;
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_clock;
//----- GPIN PORTS -----
input [0:71] gfpga_pad_RS_PREIO_A2F;
//----- GPOUT PORTS -----
output [0:71] gfpga_pad_RS_PREIO_F2A;
//----- GPOUT PORTS -----
output [0:71] gfpga_pad_RS_PREIO_SOC_CLK;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_14__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_15__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_16__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_17__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_18__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_19__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_20__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_21__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_22__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_23__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_24__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_25__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_26__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_27__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_28__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_29__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_30__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_31__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_32__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_33__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_34__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_35__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_36__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_37__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_38__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_39__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_40__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_41__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_42__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_43__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_44__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_45__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_46__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_47__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_48__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_49__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_50__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_51__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_52__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_53__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_54__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_55__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_56__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_57__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_58__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_59__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_60__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_61__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_62__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_63__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_64__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_65__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_66__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_67__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_68__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_69__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_70__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_71__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_1__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_2__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_3__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_4__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_5__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_6__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_7__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_8__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_9__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_10__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_11__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_12__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_13__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_1__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_1__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_1__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_1__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_1__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_1__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_1__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_1__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_1__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_1__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_1__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_1__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_1__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_1__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_1__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_1__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_2__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_2__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_2__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_2__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_2__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_2__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_2__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_2__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_2__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_2__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_2__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_2__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_2__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_2__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_2__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_2__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_3__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_3__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_3__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_3__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_3__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_3__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_3__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_3__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_3__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_3__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_3__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_3__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_3__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_3__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_3__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_3__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_4__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_4__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_4__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_4__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_4__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_4__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_4__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_4__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_4__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_4__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_4__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_4__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_4__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_4__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_4__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_4__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_5__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_5__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_5__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_5__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_5__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_5__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_5__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_5__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_5__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_5__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_5__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_5__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_5__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_5__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_5__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_5__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_6__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_6__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_6__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_6__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_6__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_6__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_6__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_6__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_6__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_6__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_6__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_6__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_6__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_6__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_6__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_6__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_7__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_7__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_7__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_7__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_7__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_7__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_7__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_7__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_7__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_7__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_7__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_7__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_7__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_7__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_7__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_7__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_8__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_8__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_8__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_8__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_8__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_8__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_8__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_8__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_8__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_8__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_8__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_8__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_8__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_8__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_8__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_8__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_9__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_9__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_9__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_9__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_9__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_9__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_9__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_9__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_9__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_9__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_9__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_9__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_9__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_9__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_9__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_9__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_10__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_10__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_10__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_10__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_10__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_10__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_10__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_10__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_10__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_10__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_10__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_10__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_10__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_10__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_10__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_10__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_11__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_11__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_11__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_11__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_11__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_11__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_11__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_11__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_11__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_11__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_11__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_11__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_11__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_11__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_11__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_11__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_12__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_12__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_12__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_12__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_12__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_12__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_12__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_12__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_12__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_12__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_12__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_12__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_12__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_12__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_12__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_12__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_13__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_13__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_13__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_13__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_13__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_13__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_13__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_13__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_13__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_13__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_13__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_13__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_13__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_13__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_13__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_13__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_14__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_14__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_14__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_14__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_14__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_14__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_14__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_14__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_14__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_14__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_14__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_14__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_14__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_14__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_14__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_14__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_15__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_15__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_15__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_15__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_15__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_15__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_15__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_15__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_15__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_15__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_15__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_15__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_15__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_15__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_15__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_15__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_16__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_16__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_16__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_16__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_16__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_16__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_16__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_16__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_16__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_16__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_16__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_16__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_16__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_16__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_16__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_16__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_17__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_17__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_17__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_17__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_17__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_17__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_17__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_17__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_17__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_17__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_17__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_17__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_17__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_17__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_17__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_17__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_18__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_18__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_18__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_18__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_18__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_18__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_18__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_18__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_18__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_18__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_18__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_18__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_18__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_18__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_18__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_18__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_19__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_19__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_19__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_19__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_19__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_19__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_19__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_19__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_19__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_19__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_19__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_19__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_19__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_19__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_19__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_19__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_20__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_20__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_20__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_20__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_20__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_20__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_20__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_20__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_20__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_20__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_20__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_20__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_20__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_20__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_20__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_20__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_21__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_21__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_21__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_21__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_21__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_21__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_21__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_21__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_21__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_21__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_21__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_21__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_21__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_21__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_21__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_21__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_22__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_22__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_22__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_22__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_22__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_22__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_22__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_22__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_22__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_22__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_22__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_22__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_22__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_22__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_22__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_22__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_23__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_23__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_23__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_23__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_23__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_23__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_23__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_23__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_23__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_23__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_23__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_23__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_23__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_23__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_23__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_23__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_24__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_24__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_24__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_24__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_24__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_24__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_24__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_24__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_24__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_24__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_24__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_24__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_24__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_24__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_24__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_24__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_25__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_25__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_25__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_25__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_25__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_25__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_25__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_25__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_25__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_25__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_25__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_25__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_25__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_25__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_25__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_25__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_26__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_26__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_26__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_26__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_26__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_26__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_26__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_26__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_26__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_26__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_26__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_26__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_26__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_26__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_26__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_26__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_27__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_27__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_27__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_27__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_27__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_27__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_27__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_27__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_27__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_27__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_27__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_27__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_27__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_27__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_27__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_27__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_28__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_28__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_28__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_28__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_28__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_28__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_28__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_28__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_28__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_28__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_28__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_28__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_28__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_28__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_28__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_28__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_29__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_29__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_29__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_29__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_29__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_29__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_29__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_29__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_29__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_29__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_29__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_29__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_29__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_29__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_29__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_29__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_30__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_30__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_30__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_30__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_30__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_30__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_30__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_30__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_30__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_30__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_30__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_30__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_30__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_30__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_30__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_30__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_31__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_31__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_31__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_31__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_31__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_31__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_31__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_31__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_31__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_31__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_31__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_31__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_31__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_31__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_31__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_31__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_32__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_32__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_32__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_32__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_32__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_32__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_32__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_32__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_32__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_32__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_32__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_32__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_32__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_32__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_32__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_32__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_33__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_33__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_33__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_33__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_33__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_33__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_33__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_33__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_33__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_33__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_33__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_33__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_33__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_33__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_33__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_33__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_34__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_34__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_34__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_34__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_34__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_34__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_34__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_34__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_34__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_34__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_34__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_34__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_34__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_34__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_34__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_34__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_35__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_35__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_35__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_35__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_35__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_35__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_35__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_35__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_35__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_35__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_35__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_35__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_35__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_35__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_35__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_35__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_36__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_36__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_36__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_36__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_36__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_36__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_36__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_36__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_36__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_36__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_36__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_36__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_36__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_36__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_36__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_36__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_37__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_37__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_37__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_37__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_37__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_37__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_37__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_37__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_37__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_37__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_37__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_37__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_37__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_37__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_37__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_37__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_38__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_38__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_38__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_38__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_38__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_38__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_38__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_38__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_38__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_38__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_38__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_38__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_38__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_38__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_38__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_38__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_39__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_39__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_39__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_39__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_39__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_39__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_39__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_39__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_39__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_39__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_39__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_39__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_39__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_39__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_39__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_39__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_40__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_40__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_40__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_40__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_40__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_40__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_40__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_40__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_40__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_40__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_40__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_40__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_40__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_40__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_40__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_40__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_41__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_41__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_41__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_41__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_41__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_41__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_41__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_41__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_41__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_41__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_41__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_41__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_41__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_41__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_41__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_41__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_42__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_42__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_42__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_42__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_42__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_42__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_42__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_42__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_42__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_42__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_42__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_42__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_42__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_42__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_42__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_42__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_43__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_43__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_43__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_43__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_43__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_43__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_43__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_43__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_43__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_43__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_43__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_43__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_43__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_43__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_43__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_43__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_44__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_44__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_44__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_44__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_44__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_44__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_44__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_44__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_44__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_44__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_44__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_44__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_44__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_44__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_44__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_44__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_45__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_45__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_45__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_45__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_45__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_45__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_45__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_45__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_45__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_45__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_45__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_45__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_45__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_45__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_45__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_45__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_46__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_46__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_46__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_46__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_46__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_46__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_46__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_46__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_46__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_46__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_46__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_46__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_46__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_46__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_46__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_46__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_47__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_47__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_47__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_47__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_47__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_47__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_47__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_47__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_47__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_47__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_47__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_47__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_47__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_47__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_47__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_47__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_48__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_48__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_48__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_48__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_48__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_48__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_48__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_48__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_48__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_48__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_48__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_48__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_48__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_48__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_48__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_48__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_49__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_49__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_49__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_49__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_49__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_49__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_49__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_49__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_49__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_49__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_49__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_49__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_49__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_49__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_49__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_49__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_50__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_50__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_50__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_50__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_50__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_50__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_50__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_50__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_50__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_50__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_50__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_50__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_50__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_50__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_50__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_50__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_51__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_51__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_51__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_51__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_51__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_51__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_51__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_51__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_51__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_51__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_51__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_51__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_51__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_51__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_51__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_51__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_52__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_52__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_52__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_52__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_52__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_52__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_52__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_52__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_52__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_52__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_52__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_52__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_52__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_52__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_52__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_52__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_53__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_53__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_53__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_53__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_53__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_53__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_53__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_53__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_53__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_53__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_53__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_53__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_53__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_53__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_53__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_53__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_54__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_54__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_54__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_54__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_54__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_54__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_54__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_54__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_54__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_54__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_54__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_54__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_54__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_54__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_54__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_54__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_55__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_55__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_55__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_55__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_55__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_55__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_55__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_55__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_55__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_55__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_55__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_55__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_55__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_55__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_55__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_55__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_56__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_56__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_56__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_56__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_56__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_56__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_56__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_56__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_56__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_56__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_56__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_56__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_56__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_56__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_56__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_56__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_57__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_57__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_57__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_57__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_57__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_57__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_57__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_57__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_57__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_57__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_57__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_57__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_57__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_57__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_57__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_57__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_58__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_58__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_58__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_58__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_58__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_58__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_58__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_58__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_58__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_58__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_58__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_58__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_58__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_58__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_58__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_58__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_59__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_59__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_59__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_59__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_59__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_59__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_59__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_59__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_59__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_59__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_59__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_59__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_59__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_59__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_59__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_59__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_60__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_60__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_60__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_60__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_60__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_60__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_60__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_60__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_60__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_60__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_60__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_60__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_60__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_60__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_60__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_60__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_61__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_61__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_61__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_61__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_61__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_61__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_61__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_61__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_61__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_61__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_61__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_61__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_61__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_61__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_61__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_61__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_62__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_62__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_62__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_62__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_62__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_62__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_62__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_62__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_62__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_62__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_62__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_62__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_62__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_62__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_62__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_62__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_63__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_63__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_63__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_63__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_63__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_63__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_63__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_63__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_63__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_63__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_63__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_63__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_63__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_63__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_63__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_63__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_64__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_64__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_64__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_64__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_64__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_64__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_64__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_64__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_64__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_64__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_64__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_64__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_64__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_64__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_64__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_64__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_65__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_65__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_65__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_65__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_65__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_65__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_65__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_65__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_65__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_65__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_65__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_65__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_65__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_65__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_65__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_65__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_66__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_66__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_66__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_66__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_66__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_66__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_66__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_66__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_66__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_66__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_66__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_66__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_66__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_66__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_66__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_66__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_67__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_67__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_67__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_67__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_67__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_67__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_67__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_67__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_67__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_67__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_67__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_67__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_67__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_67__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_67__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_67__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_68__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_68__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_68__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_68__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_68__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_68__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_68__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_68__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_68__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_68__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_68__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_68__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_68__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_68__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_68__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_68__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_69__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_69__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_69__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_69__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_69__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_69__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_69__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_69__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_69__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_69__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_69__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_69__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_69__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_69__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_69__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_69__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_70__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_70__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_70__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_70__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_70__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_70__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_70__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_70__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_70__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_70__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_70__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_70__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_70__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_70__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_70__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_70__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_71__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_71__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_71__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_71__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_71__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_71__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_71__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_71__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_71__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_71__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_71__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_71__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_71__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_71__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_71__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_71__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_1__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_2__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_3__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_4__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_5__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_6__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_7__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_8__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_9__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_10__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_11__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_12__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_13__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_14__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_15__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_16__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_17__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_18__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_19__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_20__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_21__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_22__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_23__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_24__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_25__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_26__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_27__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_28__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_29__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_30__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_31__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_32__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_33__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_34__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_35__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_36__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_37__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_38__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_39__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_40__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_41__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_42__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_43__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_44__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_45__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_46__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_47__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_48__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_49__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_50__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_51__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_52__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_53__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_54__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_55__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_56__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_57__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_58__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_59__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_60__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_61__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_62__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_63__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_64__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_65__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_66__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_67__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_68__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_69__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_70__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_71__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_12__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_13__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_14__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_15__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_16__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_17__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_18__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_19__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_20__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_21__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_22__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_23__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_1__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_2__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_3__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_4__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_5__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_6__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_7__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_8__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_9__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_10__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_11__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_24__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_25__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_26__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_27__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_28__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_29__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_30__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_31__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_32__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_33__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_34__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_35__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_36__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_37__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_38__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_39__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_40__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_41__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_42__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_43__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_44__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_45__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_46__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_47__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_48__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_49__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_50__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_51__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_52__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_53__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_54__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_55__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_56__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_57__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_58__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_59__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_60__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_61__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_62__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_63__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_64__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_65__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_66__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_67__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_68__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_69__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_70__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_71__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_1__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_2__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_3__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_4__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_5__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_6__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_7__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_8__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_9__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_10__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_11__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_12__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_13__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_14__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_15__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_16__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_17__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_18__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_19__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_20__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_21__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_22__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_23__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_24__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_25__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_26__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_27__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_28__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_29__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_30__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_31__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_32__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_33__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_34__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_35__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_36__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_37__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_38__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_39__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_40__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_41__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_42__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_43__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_44__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_45__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_46__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_47__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_48__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_49__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_50__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_51__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_52__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_53__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_54__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_55__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_56__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_57__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_58__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_59__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_60__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_61__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_62__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_63__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_64__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_65__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_66__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_67__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_68__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_69__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_70__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_71__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	logical_tile_io_mode_io_ logical_tile_io_mode_io__0 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[0]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[0]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[0]),
		.io_f2a_i(right_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_0__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_0__pin_clk_0_, bottom_width_0_height_0_subtile_0__pin_clk_1_, bottom_width_0_height_0_subtile_0__pin_clk_2_, bottom_width_0_height_0_subtile_0__pin_clk_3_, bottom_width_0_height_0_subtile_0__pin_clk_4_, bottom_width_0_height_0_subtile_0__pin_clk_5_, bottom_width_0_height_0_subtile_0__pin_clk_6_, bottom_width_0_height_0_subtile_0__pin_clk_7_, bottom_width_0_height_0_subtile_0__pin_clk_8_, bottom_width_0_height_0_subtile_0__pin_clk_9_, bottom_width_0_height_0_subtile_0__pin_clk_10_, bottom_width_0_height_0_subtile_0__pin_clk_11_, bottom_width_0_height_0_subtile_0__pin_clk_12_, bottom_width_0_height_0_subtile_0__pin_clk_13_, bottom_width_0_height_0_subtile_0__pin_clk_14_, bottom_width_0_height_0_subtile_0__pin_clk_15_}),
		.ccff_head(ccff_head),
		.io_a2f_o(bottom_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_0__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__0_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__1 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[1]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[1]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[1]),
		.io_f2a_i(right_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_1__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_1__pin_clk_0_, bottom_width_0_height_0_subtile_1__pin_clk_1_, bottom_width_0_height_0_subtile_1__pin_clk_2_, bottom_width_0_height_0_subtile_1__pin_clk_3_, bottom_width_0_height_0_subtile_1__pin_clk_4_, bottom_width_0_height_0_subtile_1__pin_clk_5_, bottom_width_0_height_0_subtile_1__pin_clk_6_, bottom_width_0_height_0_subtile_1__pin_clk_7_, bottom_width_0_height_0_subtile_1__pin_clk_8_, bottom_width_0_height_0_subtile_1__pin_clk_9_, bottom_width_0_height_0_subtile_1__pin_clk_10_, bottom_width_0_height_0_subtile_1__pin_clk_11_, bottom_width_0_height_0_subtile_1__pin_clk_12_, bottom_width_0_height_0_subtile_1__pin_clk_13_, bottom_width_0_height_0_subtile_1__pin_clk_14_, bottom_width_0_height_0_subtile_1__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__0_ccff_tail),
		.io_a2f_o(bottom_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_1__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__1_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__2 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[2]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[2]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[2]),
		.io_f2a_i(right_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_2__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_2__pin_clk_0_, bottom_width_0_height_0_subtile_2__pin_clk_1_, bottom_width_0_height_0_subtile_2__pin_clk_2_, bottom_width_0_height_0_subtile_2__pin_clk_3_, bottom_width_0_height_0_subtile_2__pin_clk_4_, bottom_width_0_height_0_subtile_2__pin_clk_5_, bottom_width_0_height_0_subtile_2__pin_clk_6_, bottom_width_0_height_0_subtile_2__pin_clk_7_, bottom_width_0_height_0_subtile_2__pin_clk_8_, bottom_width_0_height_0_subtile_2__pin_clk_9_, bottom_width_0_height_0_subtile_2__pin_clk_10_, bottom_width_0_height_0_subtile_2__pin_clk_11_, bottom_width_0_height_0_subtile_2__pin_clk_12_, bottom_width_0_height_0_subtile_2__pin_clk_13_, bottom_width_0_height_0_subtile_2__pin_clk_14_, bottom_width_0_height_0_subtile_2__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__1_ccff_tail),
		.io_a2f_o(bottom_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_2__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__2_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__3 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[3]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[3]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[3]),
		.io_f2a_i(right_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_3__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_3__pin_clk_0_, bottom_width_0_height_0_subtile_3__pin_clk_1_, bottom_width_0_height_0_subtile_3__pin_clk_2_, bottom_width_0_height_0_subtile_3__pin_clk_3_, bottom_width_0_height_0_subtile_3__pin_clk_4_, bottom_width_0_height_0_subtile_3__pin_clk_5_, bottom_width_0_height_0_subtile_3__pin_clk_6_, bottom_width_0_height_0_subtile_3__pin_clk_7_, bottom_width_0_height_0_subtile_3__pin_clk_8_, bottom_width_0_height_0_subtile_3__pin_clk_9_, bottom_width_0_height_0_subtile_3__pin_clk_10_, bottom_width_0_height_0_subtile_3__pin_clk_11_, bottom_width_0_height_0_subtile_3__pin_clk_12_, bottom_width_0_height_0_subtile_3__pin_clk_13_, bottom_width_0_height_0_subtile_3__pin_clk_14_, bottom_width_0_height_0_subtile_3__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__2_ccff_tail),
		.io_a2f_o(bottom_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_3__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__3_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__4 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[4]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[4]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[4]),
		.io_f2a_i(right_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_4__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_4__pin_clk_0_, bottom_width_0_height_0_subtile_4__pin_clk_1_, bottom_width_0_height_0_subtile_4__pin_clk_2_, bottom_width_0_height_0_subtile_4__pin_clk_3_, bottom_width_0_height_0_subtile_4__pin_clk_4_, bottom_width_0_height_0_subtile_4__pin_clk_5_, bottom_width_0_height_0_subtile_4__pin_clk_6_, bottom_width_0_height_0_subtile_4__pin_clk_7_, bottom_width_0_height_0_subtile_4__pin_clk_8_, bottom_width_0_height_0_subtile_4__pin_clk_9_, bottom_width_0_height_0_subtile_4__pin_clk_10_, bottom_width_0_height_0_subtile_4__pin_clk_11_, bottom_width_0_height_0_subtile_4__pin_clk_12_, bottom_width_0_height_0_subtile_4__pin_clk_13_, bottom_width_0_height_0_subtile_4__pin_clk_14_, bottom_width_0_height_0_subtile_4__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__3_ccff_tail),
		.io_a2f_o(bottom_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_4__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__4_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__5 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[5]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[5]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[5]),
		.io_f2a_i(right_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_5__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_5__pin_clk_0_, bottom_width_0_height_0_subtile_5__pin_clk_1_, bottom_width_0_height_0_subtile_5__pin_clk_2_, bottom_width_0_height_0_subtile_5__pin_clk_3_, bottom_width_0_height_0_subtile_5__pin_clk_4_, bottom_width_0_height_0_subtile_5__pin_clk_5_, bottom_width_0_height_0_subtile_5__pin_clk_6_, bottom_width_0_height_0_subtile_5__pin_clk_7_, bottom_width_0_height_0_subtile_5__pin_clk_8_, bottom_width_0_height_0_subtile_5__pin_clk_9_, bottom_width_0_height_0_subtile_5__pin_clk_10_, bottom_width_0_height_0_subtile_5__pin_clk_11_, bottom_width_0_height_0_subtile_5__pin_clk_12_, bottom_width_0_height_0_subtile_5__pin_clk_13_, bottom_width_0_height_0_subtile_5__pin_clk_14_, bottom_width_0_height_0_subtile_5__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__4_ccff_tail),
		.io_a2f_o(bottom_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_5__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__5_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__6 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[6]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[6]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[6]),
		.io_f2a_i(right_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_6__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_6__pin_clk_0_, bottom_width_0_height_0_subtile_6__pin_clk_1_, bottom_width_0_height_0_subtile_6__pin_clk_2_, bottom_width_0_height_0_subtile_6__pin_clk_3_, bottom_width_0_height_0_subtile_6__pin_clk_4_, bottom_width_0_height_0_subtile_6__pin_clk_5_, bottom_width_0_height_0_subtile_6__pin_clk_6_, bottom_width_0_height_0_subtile_6__pin_clk_7_, bottom_width_0_height_0_subtile_6__pin_clk_8_, bottom_width_0_height_0_subtile_6__pin_clk_9_, bottom_width_0_height_0_subtile_6__pin_clk_10_, bottom_width_0_height_0_subtile_6__pin_clk_11_, bottom_width_0_height_0_subtile_6__pin_clk_12_, bottom_width_0_height_0_subtile_6__pin_clk_13_, bottom_width_0_height_0_subtile_6__pin_clk_14_, bottom_width_0_height_0_subtile_6__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__5_ccff_tail),
		.io_a2f_o(bottom_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_6__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__6_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__7 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[7]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[7]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[7]),
		.io_f2a_i(right_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_7__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_7__pin_clk_0_, bottom_width_0_height_0_subtile_7__pin_clk_1_, bottom_width_0_height_0_subtile_7__pin_clk_2_, bottom_width_0_height_0_subtile_7__pin_clk_3_, bottom_width_0_height_0_subtile_7__pin_clk_4_, bottom_width_0_height_0_subtile_7__pin_clk_5_, bottom_width_0_height_0_subtile_7__pin_clk_6_, bottom_width_0_height_0_subtile_7__pin_clk_7_, bottom_width_0_height_0_subtile_7__pin_clk_8_, bottom_width_0_height_0_subtile_7__pin_clk_9_, bottom_width_0_height_0_subtile_7__pin_clk_10_, bottom_width_0_height_0_subtile_7__pin_clk_11_, bottom_width_0_height_0_subtile_7__pin_clk_12_, bottom_width_0_height_0_subtile_7__pin_clk_13_, bottom_width_0_height_0_subtile_7__pin_clk_14_, bottom_width_0_height_0_subtile_7__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__6_ccff_tail),
		.io_a2f_o(bottom_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_7__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__7_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__8 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[8]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[8]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[8]),
		.io_f2a_i(right_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_8__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_8__pin_clk_0_, bottom_width_0_height_0_subtile_8__pin_clk_1_, bottom_width_0_height_0_subtile_8__pin_clk_2_, bottom_width_0_height_0_subtile_8__pin_clk_3_, bottom_width_0_height_0_subtile_8__pin_clk_4_, bottom_width_0_height_0_subtile_8__pin_clk_5_, bottom_width_0_height_0_subtile_8__pin_clk_6_, bottom_width_0_height_0_subtile_8__pin_clk_7_, bottom_width_0_height_0_subtile_8__pin_clk_8_, bottom_width_0_height_0_subtile_8__pin_clk_9_, bottom_width_0_height_0_subtile_8__pin_clk_10_, bottom_width_0_height_0_subtile_8__pin_clk_11_, bottom_width_0_height_0_subtile_8__pin_clk_12_, bottom_width_0_height_0_subtile_8__pin_clk_13_, bottom_width_0_height_0_subtile_8__pin_clk_14_, bottom_width_0_height_0_subtile_8__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__7_ccff_tail),
		.io_a2f_o(bottom_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_8__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__8_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__9 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[9]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[9]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[9]),
		.io_f2a_i(right_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_9__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_9__pin_clk_0_, bottom_width_0_height_0_subtile_9__pin_clk_1_, bottom_width_0_height_0_subtile_9__pin_clk_2_, bottom_width_0_height_0_subtile_9__pin_clk_3_, bottom_width_0_height_0_subtile_9__pin_clk_4_, bottom_width_0_height_0_subtile_9__pin_clk_5_, bottom_width_0_height_0_subtile_9__pin_clk_6_, bottom_width_0_height_0_subtile_9__pin_clk_7_, bottom_width_0_height_0_subtile_9__pin_clk_8_, bottom_width_0_height_0_subtile_9__pin_clk_9_, bottom_width_0_height_0_subtile_9__pin_clk_10_, bottom_width_0_height_0_subtile_9__pin_clk_11_, bottom_width_0_height_0_subtile_9__pin_clk_12_, bottom_width_0_height_0_subtile_9__pin_clk_13_, bottom_width_0_height_0_subtile_9__pin_clk_14_, bottom_width_0_height_0_subtile_9__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__8_ccff_tail),
		.io_a2f_o(bottom_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_9__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__9_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__10 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[10]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[10]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[10]),
		.io_f2a_i(right_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_10__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_10__pin_clk_0_, bottom_width_0_height_0_subtile_10__pin_clk_1_, bottom_width_0_height_0_subtile_10__pin_clk_2_, bottom_width_0_height_0_subtile_10__pin_clk_3_, bottom_width_0_height_0_subtile_10__pin_clk_4_, bottom_width_0_height_0_subtile_10__pin_clk_5_, bottom_width_0_height_0_subtile_10__pin_clk_6_, bottom_width_0_height_0_subtile_10__pin_clk_7_, bottom_width_0_height_0_subtile_10__pin_clk_8_, bottom_width_0_height_0_subtile_10__pin_clk_9_, bottom_width_0_height_0_subtile_10__pin_clk_10_, bottom_width_0_height_0_subtile_10__pin_clk_11_, bottom_width_0_height_0_subtile_10__pin_clk_12_, bottom_width_0_height_0_subtile_10__pin_clk_13_, bottom_width_0_height_0_subtile_10__pin_clk_14_, bottom_width_0_height_0_subtile_10__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__9_ccff_tail),
		.io_a2f_o(bottom_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_10__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__10_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__11 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[11]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[11]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[11]),
		.io_f2a_i(right_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_11__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_11__pin_clk_0_, bottom_width_0_height_0_subtile_11__pin_clk_1_, bottom_width_0_height_0_subtile_11__pin_clk_2_, bottom_width_0_height_0_subtile_11__pin_clk_3_, bottom_width_0_height_0_subtile_11__pin_clk_4_, bottom_width_0_height_0_subtile_11__pin_clk_5_, bottom_width_0_height_0_subtile_11__pin_clk_6_, bottom_width_0_height_0_subtile_11__pin_clk_7_, bottom_width_0_height_0_subtile_11__pin_clk_8_, bottom_width_0_height_0_subtile_11__pin_clk_9_, bottom_width_0_height_0_subtile_11__pin_clk_10_, bottom_width_0_height_0_subtile_11__pin_clk_11_, bottom_width_0_height_0_subtile_11__pin_clk_12_, bottom_width_0_height_0_subtile_11__pin_clk_13_, bottom_width_0_height_0_subtile_11__pin_clk_14_, bottom_width_0_height_0_subtile_11__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__10_ccff_tail),
		.io_a2f_o(bottom_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_11__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__11_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__12 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[12]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[12]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[12]),
		.io_f2a_i(right_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_12__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_12__pin_clk_0_, bottom_width_0_height_0_subtile_12__pin_clk_1_, bottom_width_0_height_0_subtile_12__pin_clk_2_, bottom_width_0_height_0_subtile_12__pin_clk_3_, bottom_width_0_height_0_subtile_12__pin_clk_4_, bottom_width_0_height_0_subtile_12__pin_clk_5_, bottom_width_0_height_0_subtile_12__pin_clk_6_, bottom_width_0_height_0_subtile_12__pin_clk_7_, bottom_width_0_height_0_subtile_12__pin_clk_8_, bottom_width_0_height_0_subtile_12__pin_clk_9_, bottom_width_0_height_0_subtile_12__pin_clk_10_, bottom_width_0_height_0_subtile_12__pin_clk_11_, bottom_width_0_height_0_subtile_12__pin_clk_12_, bottom_width_0_height_0_subtile_12__pin_clk_13_, bottom_width_0_height_0_subtile_12__pin_clk_14_, bottom_width_0_height_0_subtile_12__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__11_ccff_tail),
		.io_a2f_o(right_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_12__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__12_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__13 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[13]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[13]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[13]),
		.io_f2a_i(right_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_13__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_13__pin_clk_0_, bottom_width_0_height_0_subtile_13__pin_clk_1_, bottom_width_0_height_0_subtile_13__pin_clk_2_, bottom_width_0_height_0_subtile_13__pin_clk_3_, bottom_width_0_height_0_subtile_13__pin_clk_4_, bottom_width_0_height_0_subtile_13__pin_clk_5_, bottom_width_0_height_0_subtile_13__pin_clk_6_, bottom_width_0_height_0_subtile_13__pin_clk_7_, bottom_width_0_height_0_subtile_13__pin_clk_8_, bottom_width_0_height_0_subtile_13__pin_clk_9_, bottom_width_0_height_0_subtile_13__pin_clk_10_, bottom_width_0_height_0_subtile_13__pin_clk_11_, bottom_width_0_height_0_subtile_13__pin_clk_12_, bottom_width_0_height_0_subtile_13__pin_clk_13_, bottom_width_0_height_0_subtile_13__pin_clk_14_, bottom_width_0_height_0_subtile_13__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__12_ccff_tail),
		.io_a2f_o(right_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_13__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__13_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__14 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[14]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[14]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[14]),
		.io_f2a_i(top_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_14__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_14__pin_clk_0_, bottom_width_0_height_0_subtile_14__pin_clk_1_, bottom_width_0_height_0_subtile_14__pin_clk_2_, bottom_width_0_height_0_subtile_14__pin_clk_3_, bottom_width_0_height_0_subtile_14__pin_clk_4_, bottom_width_0_height_0_subtile_14__pin_clk_5_, bottom_width_0_height_0_subtile_14__pin_clk_6_, bottom_width_0_height_0_subtile_14__pin_clk_7_, bottom_width_0_height_0_subtile_14__pin_clk_8_, bottom_width_0_height_0_subtile_14__pin_clk_9_, bottom_width_0_height_0_subtile_14__pin_clk_10_, bottom_width_0_height_0_subtile_14__pin_clk_11_, bottom_width_0_height_0_subtile_14__pin_clk_12_, bottom_width_0_height_0_subtile_14__pin_clk_13_, bottom_width_0_height_0_subtile_14__pin_clk_14_, bottom_width_0_height_0_subtile_14__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__13_ccff_tail),
		.io_a2f_o(right_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_14__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__14_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__15 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[15]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[15]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[15]),
		.io_f2a_i(top_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_15__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_15__pin_clk_0_, bottom_width_0_height_0_subtile_15__pin_clk_1_, bottom_width_0_height_0_subtile_15__pin_clk_2_, bottom_width_0_height_0_subtile_15__pin_clk_3_, bottom_width_0_height_0_subtile_15__pin_clk_4_, bottom_width_0_height_0_subtile_15__pin_clk_5_, bottom_width_0_height_0_subtile_15__pin_clk_6_, bottom_width_0_height_0_subtile_15__pin_clk_7_, bottom_width_0_height_0_subtile_15__pin_clk_8_, bottom_width_0_height_0_subtile_15__pin_clk_9_, bottom_width_0_height_0_subtile_15__pin_clk_10_, bottom_width_0_height_0_subtile_15__pin_clk_11_, bottom_width_0_height_0_subtile_15__pin_clk_12_, bottom_width_0_height_0_subtile_15__pin_clk_13_, bottom_width_0_height_0_subtile_15__pin_clk_14_, bottom_width_0_height_0_subtile_15__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__14_ccff_tail),
		.io_a2f_o(right_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_15__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__15_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__16 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[16]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[16]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[16]),
		.io_f2a_i(top_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_16__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_16__pin_clk_0_, bottom_width_0_height_0_subtile_16__pin_clk_1_, bottom_width_0_height_0_subtile_16__pin_clk_2_, bottom_width_0_height_0_subtile_16__pin_clk_3_, bottom_width_0_height_0_subtile_16__pin_clk_4_, bottom_width_0_height_0_subtile_16__pin_clk_5_, bottom_width_0_height_0_subtile_16__pin_clk_6_, bottom_width_0_height_0_subtile_16__pin_clk_7_, bottom_width_0_height_0_subtile_16__pin_clk_8_, bottom_width_0_height_0_subtile_16__pin_clk_9_, bottom_width_0_height_0_subtile_16__pin_clk_10_, bottom_width_0_height_0_subtile_16__pin_clk_11_, bottom_width_0_height_0_subtile_16__pin_clk_12_, bottom_width_0_height_0_subtile_16__pin_clk_13_, bottom_width_0_height_0_subtile_16__pin_clk_14_, bottom_width_0_height_0_subtile_16__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__15_ccff_tail),
		.io_a2f_o(right_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_16__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__16_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__17 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[17]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[17]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[17]),
		.io_f2a_i(top_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_17__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_17__pin_clk_0_, bottom_width_0_height_0_subtile_17__pin_clk_1_, bottom_width_0_height_0_subtile_17__pin_clk_2_, bottom_width_0_height_0_subtile_17__pin_clk_3_, bottom_width_0_height_0_subtile_17__pin_clk_4_, bottom_width_0_height_0_subtile_17__pin_clk_5_, bottom_width_0_height_0_subtile_17__pin_clk_6_, bottom_width_0_height_0_subtile_17__pin_clk_7_, bottom_width_0_height_0_subtile_17__pin_clk_8_, bottom_width_0_height_0_subtile_17__pin_clk_9_, bottom_width_0_height_0_subtile_17__pin_clk_10_, bottom_width_0_height_0_subtile_17__pin_clk_11_, bottom_width_0_height_0_subtile_17__pin_clk_12_, bottom_width_0_height_0_subtile_17__pin_clk_13_, bottom_width_0_height_0_subtile_17__pin_clk_14_, bottom_width_0_height_0_subtile_17__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__16_ccff_tail),
		.io_a2f_o(right_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_17__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__17_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__18 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[18]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[18]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[18]),
		.io_f2a_i(top_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_18__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_18__pin_clk_0_, bottom_width_0_height_0_subtile_18__pin_clk_1_, bottom_width_0_height_0_subtile_18__pin_clk_2_, bottom_width_0_height_0_subtile_18__pin_clk_3_, bottom_width_0_height_0_subtile_18__pin_clk_4_, bottom_width_0_height_0_subtile_18__pin_clk_5_, bottom_width_0_height_0_subtile_18__pin_clk_6_, bottom_width_0_height_0_subtile_18__pin_clk_7_, bottom_width_0_height_0_subtile_18__pin_clk_8_, bottom_width_0_height_0_subtile_18__pin_clk_9_, bottom_width_0_height_0_subtile_18__pin_clk_10_, bottom_width_0_height_0_subtile_18__pin_clk_11_, bottom_width_0_height_0_subtile_18__pin_clk_12_, bottom_width_0_height_0_subtile_18__pin_clk_13_, bottom_width_0_height_0_subtile_18__pin_clk_14_, bottom_width_0_height_0_subtile_18__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__17_ccff_tail),
		.io_a2f_o(right_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_18__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__18_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__19 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[19]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[19]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[19]),
		.io_f2a_i(top_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_19__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_19__pin_clk_0_, bottom_width_0_height_0_subtile_19__pin_clk_1_, bottom_width_0_height_0_subtile_19__pin_clk_2_, bottom_width_0_height_0_subtile_19__pin_clk_3_, bottom_width_0_height_0_subtile_19__pin_clk_4_, bottom_width_0_height_0_subtile_19__pin_clk_5_, bottom_width_0_height_0_subtile_19__pin_clk_6_, bottom_width_0_height_0_subtile_19__pin_clk_7_, bottom_width_0_height_0_subtile_19__pin_clk_8_, bottom_width_0_height_0_subtile_19__pin_clk_9_, bottom_width_0_height_0_subtile_19__pin_clk_10_, bottom_width_0_height_0_subtile_19__pin_clk_11_, bottom_width_0_height_0_subtile_19__pin_clk_12_, bottom_width_0_height_0_subtile_19__pin_clk_13_, bottom_width_0_height_0_subtile_19__pin_clk_14_, bottom_width_0_height_0_subtile_19__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__18_ccff_tail),
		.io_a2f_o(right_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_19__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__19_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__20 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[20]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[20]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[20]),
		.io_f2a_i(top_width_0_height_0_subtile_20__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_20__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_20__pin_clk_0_, bottom_width_0_height_0_subtile_20__pin_clk_1_, bottom_width_0_height_0_subtile_20__pin_clk_2_, bottom_width_0_height_0_subtile_20__pin_clk_3_, bottom_width_0_height_0_subtile_20__pin_clk_4_, bottom_width_0_height_0_subtile_20__pin_clk_5_, bottom_width_0_height_0_subtile_20__pin_clk_6_, bottom_width_0_height_0_subtile_20__pin_clk_7_, bottom_width_0_height_0_subtile_20__pin_clk_8_, bottom_width_0_height_0_subtile_20__pin_clk_9_, bottom_width_0_height_0_subtile_20__pin_clk_10_, bottom_width_0_height_0_subtile_20__pin_clk_11_, bottom_width_0_height_0_subtile_20__pin_clk_12_, bottom_width_0_height_0_subtile_20__pin_clk_13_, bottom_width_0_height_0_subtile_20__pin_clk_14_, bottom_width_0_height_0_subtile_20__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__19_ccff_tail),
		.io_a2f_o(right_width_0_height_0_subtile_20__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_20__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__20_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__21 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[21]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[21]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[21]),
		.io_f2a_i(top_width_0_height_0_subtile_21__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_21__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_21__pin_clk_0_, bottom_width_0_height_0_subtile_21__pin_clk_1_, bottom_width_0_height_0_subtile_21__pin_clk_2_, bottom_width_0_height_0_subtile_21__pin_clk_3_, bottom_width_0_height_0_subtile_21__pin_clk_4_, bottom_width_0_height_0_subtile_21__pin_clk_5_, bottom_width_0_height_0_subtile_21__pin_clk_6_, bottom_width_0_height_0_subtile_21__pin_clk_7_, bottom_width_0_height_0_subtile_21__pin_clk_8_, bottom_width_0_height_0_subtile_21__pin_clk_9_, bottom_width_0_height_0_subtile_21__pin_clk_10_, bottom_width_0_height_0_subtile_21__pin_clk_11_, bottom_width_0_height_0_subtile_21__pin_clk_12_, bottom_width_0_height_0_subtile_21__pin_clk_13_, bottom_width_0_height_0_subtile_21__pin_clk_14_, bottom_width_0_height_0_subtile_21__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__20_ccff_tail),
		.io_a2f_o(right_width_0_height_0_subtile_21__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_21__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__21_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__22 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[22]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[22]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[22]),
		.io_f2a_i(top_width_0_height_0_subtile_22__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_22__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_22__pin_clk_0_, bottom_width_0_height_0_subtile_22__pin_clk_1_, bottom_width_0_height_0_subtile_22__pin_clk_2_, bottom_width_0_height_0_subtile_22__pin_clk_3_, bottom_width_0_height_0_subtile_22__pin_clk_4_, bottom_width_0_height_0_subtile_22__pin_clk_5_, bottom_width_0_height_0_subtile_22__pin_clk_6_, bottom_width_0_height_0_subtile_22__pin_clk_7_, bottom_width_0_height_0_subtile_22__pin_clk_8_, bottom_width_0_height_0_subtile_22__pin_clk_9_, bottom_width_0_height_0_subtile_22__pin_clk_10_, bottom_width_0_height_0_subtile_22__pin_clk_11_, bottom_width_0_height_0_subtile_22__pin_clk_12_, bottom_width_0_height_0_subtile_22__pin_clk_13_, bottom_width_0_height_0_subtile_22__pin_clk_14_, bottom_width_0_height_0_subtile_22__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__21_ccff_tail),
		.io_a2f_o(right_width_0_height_0_subtile_22__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_22__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__22_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__23 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[23]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[23]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[23]),
		.io_f2a_i(top_width_0_height_0_subtile_23__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_23__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_23__pin_clk_0_, bottom_width_0_height_0_subtile_23__pin_clk_1_, bottom_width_0_height_0_subtile_23__pin_clk_2_, bottom_width_0_height_0_subtile_23__pin_clk_3_, bottom_width_0_height_0_subtile_23__pin_clk_4_, bottom_width_0_height_0_subtile_23__pin_clk_5_, bottom_width_0_height_0_subtile_23__pin_clk_6_, bottom_width_0_height_0_subtile_23__pin_clk_7_, bottom_width_0_height_0_subtile_23__pin_clk_8_, bottom_width_0_height_0_subtile_23__pin_clk_9_, bottom_width_0_height_0_subtile_23__pin_clk_10_, bottom_width_0_height_0_subtile_23__pin_clk_11_, bottom_width_0_height_0_subtile_23__pin_clk_12_, bottom_width_0_height_0_subtile_23__pin_clk_13_, bottom_width_0_height_0_subtile_23__pin_clk_14_, bottom_width_0_height_0_subtile_23__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__22_ccff_tail),
		.io_a2f_o(right_width_0_height_0_subtile_23__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_23__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__23_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__24 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[24]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[24]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[24]),
		.io_f2a_i(top_width_0_height_0_subtile_24__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_24__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_24__pin_clk_0_, bottom_width_0_height_0_subtile_24__pin_clk_1_, bottom_width_0_height_0_subtile_24__pin_clk_2_, bottom_width_0_height_0_subtile_24__pin_clk_3_, bottom_width_0_height_0_subtile_24__pin_clk_4_, bottom_width_0_height_0_subtile_24__pin_clk_5_, bottom_width_0_height_0_subtile_24__pin_clk_6_, bottom_width_0_height_0_subtile_24__pin_clk_7_, bottom_width_0_height_0_subtile_24__pin_clk_8_, bottom_width_0_height_0_subtile_24__pin_clk_9_, bottom_width_0_height_0_subtile_24__pin_clk_10_, bottom_width_0_height_0_subtile_24__pin_clk_11_, bottom_width_0_height_0_subtile_24__pin_clk_12_, bottom_width_0_height_0_subtile_24__pin_clk_13_, bottom_width_0_height_0_subtile_24__pin_clk_14_, bottom_width_0_height_0_subtile_24__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__23_ccff_tail),
		.io_a2f_o(bottom_width_0_height_0_subtile_24__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_24__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__24_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__25 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[25]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[25]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[25]),
		.io_f2a_i(top_width_0_height_0_subtile_25__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_25__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_25__pin_clk_0_, bottom_width_0_height_0_subtile_25__pin_clk_1_, bottom_width_0_height_0_subtile_25__pin_clk_2_, bottom_width_0_height_0_subtile_25__pin_clk_3_, bottom_width_0_height_0_subtile_25__pin_clk_4_, bottom_width_0_height_0_subtile_25__pin_clk_5_, bottom_width_0_height_0_subtile_25__pin_clk_6_, bottom_width_0_height_0_subtile_25__pin_clk_7_, bottom_width_0_height_0_subtile_25__pin_clk_8_, bottom_width_0_height_0_subtile_25__pin_clk_9_, bottom_width_0_height_0_subtile_25__pin_clk_10_, bottom_width_0_height_0_subtile_25__pin_clk_11_, bottom_width_0_height_0_subtile_25__pin_clk_12_, bottom_width_0_height_0_subtile_25__pin_clk_13_, bottom_width_0_height_0_subtile_25__pin_clk_14_, bottom_width_0_height_0_subtile_25__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__24_ccff_tail),
		.io_a2f_o(bottom_width_0_height_0_subtile_25__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_25__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__25_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__26 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[26]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[26]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[26]),
		.io_f2a_i(top_width_0_height_0_subtile_26__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_26__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_26__pin_clk_0_, bottom_width_0_height_0_subtile_26__pin_clk_1_, bottom_width_0_height_0_subtile_26__pin_clk_2_, bottom_width_0_height_0_subtile_26__pin_clk_3_, bottom_width_0_height_0_subtile_26__pin_clk_4_, bottom_width_0_height_0_subtile_26__pin_clk_5_, bottom_width_0_height_0_subtile_26__pin_clk_6_, bottom_width_0_height_0_subtile_26__pin_clk_7_, bottom_width_0_height_0_subtile_26__pin_clk_8_, bottom_width_0_height_0_subtile_26__pin_clk_9_, bottom_width_0_height_0_subtile_26__pin_clk_10_, bottom_width_0_height_0_subtile_26__pin_clk_11_, bottom_width_0_height_0_subtile_26__pin_clk_12_, bottom_width_0_height_0_subtile_26__pin_clk_13_, bottom_width_0_height_0_subtile_26__pin_clk_14_, bottom_width_0_height_0_subtile_26__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__25_ccff_tail),
		.io_a2f_o(bottom_width_0_height_0_subtile_26__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_26__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__26_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__27 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[27]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[27]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[27]),
		.io_f2a_i(top_width_0_height_0_subtile_27__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_27__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_27__pin_clk_0_, bottom_width_0_height_0_subtile_27__pin_clk_1_, bottom_width_0_height_0_subtile_27__pin_clk_2_, bottom_width_0_height_0_subtile_27__pin_clk_3_, bottom_width_0_height_0_subtile_27__pin_clk_4_, bottom_width_0_height_0_subtile_27__pin_clk_5_, bottom_width_0_height_0_subtile_27__pin_clk_6_, bottom_width_0_height_0_subtile_27__pin_clk_7_, bottom_width_0_height_0_subtile_27__pin_clk_8_, bottom_width_0_height_0_subtile_27__pin_clk_9_, bottom_width_0_height_0_subtile_27__pin_clk_10_, bottom_width_0_height_0_subtile_27__pin_clk_11_, bottom_width_0_height_0_subtile_27__pin_clk_12_, bottom_width_0_height_0_subtile_27__pin_clk_13_, bottom_width_0_height_0_subtile_27__pin_clk_14_, bottom_width_0_height_0_subtile_27__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__26_ccff_tail),
		.io_a2f_o(bottom_width_0_height_0_subtile_27__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_27__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__27_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__28 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[28]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[28]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[28]),
		.io_f2a_i(top_width_0_height_0_subtile_28__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_28__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_28__pin_clk_0_, bottom_width_0_height_0_subtile_28__pin_clk_1_, bottom_width_0_height_0_subtile_28__pin_clk_2_, bottom_width_0_height_0_subtile_28__pin_clk_3_, bottom_width_0_height_0_subtile_28__pin_clk_4_, bottom_width_0_height_0_subtile_28__pin_clk_5_, bottom_width_0_height_0_subtile_28__pin_clk_6_, bottom_width_0_height_0_subtile_28__pin_clk_7_, bottom_width_0_height_0_subtile_28__pin_clk_8_, bottom_width_0_height_0_subtile_28__pin_clk_9_, bottom_width_0_height_0_subtile_28__pin_clk_10_, bottom_width_0_height_0_subtile_28__pin_clk_11_, bottom_width_0_height_0_subtile_28__pin_clk_12_, bottom_width_0_height_0_subtile_28__pin_clk_13_, bottom_width_0_height_0_subtile_28__pin_clk_14_, bottom_width_0_height_0_subtile_28__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__27_ccff_tail),
		.io_a2f_o(bottom_width_0_height_0_subtile_28__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_28__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__28_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__29 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[29]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[29]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[29]),
		.io_f2a_i(top_width_0_height_0_subtile_29__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_29__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_29__pin_clk_0_, bottom_width_0_height_0_subtile_29__pin_clk_1_, bottom_width_0_height_0_subtile_29__pin_clk_2_, bottom_width_0_height_0_subtile_29__pin_clk_3_, bottom_width_0_height_0_subtile_29__pin_clk_4_, bottom_width_0_height_0_subtile_29__pin_clk_5_, bottom_width_0_height_0_subtile_29__pin_clk_6_, bottom_width_0_height_0_subtile_29__pin_clk_7_, bottom_width_0_height_0_subtile_29__pin_clk_8_, bottom_width_0_height_0_subtile_29__pin_clk_9_, bottom_width_0_height_0_subtile_29__pin_clk_10_, bottom_width_0_height_0_subtile_29__pin_clk_11_, bottom_width_0_height_0_subtile_29__pin_clk_12_, bottom_width_0_height_0_subtile_29__pin_clk_13_, bottom_width_0_height_0_subtile_29__pin_clk_14_, bottom_width_0_height_0_subtile_29__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__28_ccff_tail),
		.io_a2f_o(bottom_width_0_height_0_subtile_29__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_29__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__29_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__30 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[30]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[30]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[30]),
		.io_f2a_i(top_width_0_height_0_subtile_30__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_30__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_30__pin_clk_0_, bottom_width_0_height_0_subtile_30__pin_clk_1_, bottom_width_0_height_0_subtile_30__pin_clk_2_, bottom_width_0_height_0_subtile_30__pin_clk_3_, bottom_width_0_height_0_subtile_30__pin_clk_4_, bottom_width_0_height_0_subtile_30__pin_clk_5_, bottom_width_0_height_0_subtile_30__pin_clk_6_, bottom_width_0_height_0_subtile_30__pin_clk_7_, bottom_width_0_height_0_subtile_30__pin_clk_8_, bottom_width_0_height_0_subtile_30__pin_clk_9_, bottom_width_0_height_0_subtile_30__pin_clk_10_, bottom_width_0_height_0_subtile_30__pin_clk_11_, bottom_width_0_height_0_subtile_30__pin_clk_12_, bottom_width_0_height_0_subtile_30__pin_clk_13_, bottom_width_0_height_0_subtile_30__pin_clk_14_, bottom_width_0_height_0_subtile_30__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__29_ccff_tail),
		.io_a2f_o(bottom_width_0_height_0_subtile_30__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_30__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__30_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__31 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[31]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[31]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[31]),
		.io_f2a_i(top_width_0_height_0_subtile_31__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_31__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_31__pin_clk_0_, bottom_width_0_height_0_subtile_31__pin_clk_1_, bottom_width_0_height_0_subtile_31__pin_clk_2_, bottom_width_0_height_0_subtile_31__pin_clk_3_, bottom_width_0_height_0_subtile_31__pin_clk_4_, bottom_width_0_height_0_subtile_31__pin_clk_5_, bottom_width_0_height_0_subtile_31__pin_clk_6_, bottom_width_0_height_0_subtile_31__pin_clk_7_, bottom_width_0_height_0_subtile_31__pin_clk_8_, bottom_width_0_height_0_subtile_31__pin_clk_9_, bottom_width_0_height_0_subtile_31__pin_clk_10_, bottom_width_0_height_0_subtile_31__pin_clk_11_, bottom_width_0_height_0_subtile_31__pin_clk_12_, bottom_width_0_height_0_subtile_31__pin_clk_13_, bottom_width_0_height_0_subtile_31__pin_clk_14_, bottom_width_0_height_0_subtile_31__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__30_ccff_tail),
		.io_a2f_o(bottom_width_0_height_0_subtile_31__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_31__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__31_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__32 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[32]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[32]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[32]),
		.io_f2a_i(top_width_0_height_0_subtile_32__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_32__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_32__pin_clk_0_, bottom_width_0_height_0_subtile_32__pin_clk_1_, bottom_width_0_height_0_subtile_32__pin_clk_2_, bottom_width_0_height_0_subtile_32__pin_clk_3_, bottom_width_0_height_0_subtile_32__pin_clk_4_, bottom_width_0_height_0_subtile_32__pin_clk_5_, bottom_width_0_height_0_subtile_32__pin_clk_6_, bottom_width_0_height_0_subtile_32__pin_clk_7_, bottom_width_0_height_0_subtile_32__pin_clk_8_, bottom_width_0_height_0_subtile_32__pin_clk_9_, bottom_width_0_height_0_subtile_32__pin_clk_10_, bottom_width_0_height_0_subtile_32__pin_clk_11_, bottom_width_0_height_0_subtile_32__pin_clk_12_, bottom_width_0_height_0_subtile_32__pin_clk_13_, bottom_width_0_height_0_subtile_32__pin_clk_14_, bottom_width_0_height_0_subtile_32__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__31_ccff_tail),
		.io_a2f_o(bottom_width_0_height_0_subtile_32__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_32__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__32_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__33 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[33]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[33]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[33]),
		.io_f2a_i(top_width_0_height_0_subtile_33__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_33__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_33__pin_clk_0_, bottom_width_0_height_0_subtile_33__pin_clk_1_, bottom_width_0_height_0_subtile_33__pin_clk_2_, bottom_width_0_height_0_subtile_33__pin_clk_3_, bottom_width_0_height_0_subtile_33__pin_clk_4_, bottom_width_0_height_0_subtile_33__pin_clk_5_, bottom_width_0_height_0_subtile_33__pin_clk_6_, bottom_width_0_height_0_subtile_33__pin_clk_7_, bottom_width_0_height_0_subtile_33__pin_clk_8_, bottom_width_0_height_0_subtile_33__pin_clk_9_, bottom_width_0_height_0_subtile_33__pin_clk_10_, bottom_width_0_height_0_subtile_33__pin_clk_11_, bottom_width_0_height_0_subtile_33__pin_clk_12_, bottom_width_0_height_0_subtile_33__pin_clk_13_, bottom_width_0_height_0_subtile_33__pin_clk_14_, bottom_width_0_height_0_subtile_33__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__32_ccff_tail),
		.io_a2f_o(bottom_width_0_height_0_subtile_33__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_33__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__33_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__34 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[34]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[34]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[34]),
		.io_f2a_i(top_width_0_height_0_subtile_34__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_34__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_34__pin_clk_0_, bottom_width_0_height_0_subtile_34__pin_clk_1_, bottom_width_0_height_0_subtile_34__pin_clk_2_, bottom_width_0_height_0_subtile_34__pin_clk_3_, bottom_width_0_height_0_subtile_34__pin_clk_4_, bottom_width_0_height_0_subtile_34__pin_clk_5_, bottom_width_0_height_0_subtile_34__pin_clk_6_, bottom_width_0_height_0_subtile_34__pin_clk_7_, bottom_width_0_height_0_subtile_34__pin_clk_8_, bottom_width_0_height_0_subtile_34__pin_clk_9_, bottom_width_0_height_0_subtile_34__pin_clk_10_, bottom_width_0_height_0_subtile_34__pin_clk_11_, bottom_width_0_height_0_subtile_34__pin_clk_12_, bottom_width_0_height_0_subtile_34__pin_clk_13_, bottom_width_0_height_0_subtile_34__pin_clk_14_, bottom_width_0_height_0_subtile_34__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__33_ccff_tail),
		.io_a2f_o(bottom_width_0_height_0_subtile_34__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_34__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__34_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__35 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[35]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[35]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[35]),
		.io_f2a_i(top_width_0_height_0_subtile_35__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_35__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_35__pin_clk_0_, bottom_width_0_height_0_subtile_35__pin_clk_1_, bottom_width_0_height_0_subtile_35__pin_clk_2_, bottom_width_0_height_0_subtile_35__pin_clk_3_, bottom_width_0_height_0_subtile_35__pin_clk_4_, bottom_width_0_height_0_subtile_35__pin_clk_5_, bottom_width_0_height_0_subtile_35__pin_clk_6_, bottom_width_0_height_0_subtile_35__pin_clk_7_, bottom_width_0_height_0_subtile_35__pin_clk_8_, bottom_width_0_height_0_subtile_35__pin_clk_9_, bottom_width_0_height_0_subtile_35__pin_clk_10_, bottom_width_0_height_0_subtile_35__pin_clk_11_, bottom_width_0_height_0_subtile_35__pin_clk_12_, bottom_width_0_height_0_subtile_35__pin_clk_13_, bottom_width_0_height_0_subtile_35__pin_clk_14_, bottom_width_0_height_0_subtile_35__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__34_ccff_tail),
		.io_a2f_o(bottom_width_0_height_0_subtile_35__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_35__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__35_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__36 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[36]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[36]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[36]),
		.io_f2a_i(top_width_0_height_0_subtile_36__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_36__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_36__pin_clk_0_, bottom_width_0_height_0_subtile_36__pin_clk_1_, bottom_width_0_height_0_subtile_36__pin_clk_2_, bottom_width_0_height_0_subtile_36__pin_clk_3_, bottom_width_0_height_0_subtile_36__pin_clk_4_, bottom_width_0_height_0_subtile_36__pin_clk_5_, bottom_width_0_height_0_subtile_36__pin_clk_6_, bottom_width_0_height_0_subtile_36__pin_clk_7_, bottom_width_0_height_0_subtile_36__pin_clk_8_, bottom_width_0_height_0_subtile_36__pin_clk_9_, bottom_width_0_height_0_subtile_36__pin_clk_10_, bottom_width_0_height_0_subtile_36__pin_clk_11_, bottom_width_0_height_0_subtile_36__pin_clk_12_, bottom_width_0_height_0_subtile_36__pin_clk_13_, bottom_width_0_height_0_subtile_36__pin_clk_14_, bottom_width_0_height_0_subtile_36__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__35_ccff_tail),
		.io_a2f_o(bottom_width_0_height_0_subtile_36__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_36__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__36_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__37 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[37]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[37]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[37]),
		.io_f2a_i(top_width_0_height_0_subtile_37__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_37__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_37__pin_clk_0_, bottom_width_0_height_0_subtile_37__pin_clk_1_, bottom_width_0_height_0_subtile_37__pin_clk_2_, bottom_width_0_height_0_subtile_37__pin_clk_3_, bottom_width_0_height_0_subtile_37__pin_clk_4_, bottom_width_0_height_0_subtile_37__pin_clk_5_, bottom_width_0_height_0_subtile_37__pin_clk_6_, bottom_width_0_height_0_subtile_37__pin_clk_7_, bottom_width_0_height_0_subtile_37__pin_clk_8_, bottom_width_0_height_0_subtile_37__pin_clk_9_, bottom_width_0_height_0_subtile_37__pin_clk_10_, bottom_width_0_height_0_subtile_37__pin_clk_11_, bottom_width_0_height_0_subtile_37__pin_clk_12_, bottom_width_0_height_0_subtile_37__pin_clk_13_, bottom_width_0_height_0_subtile_37__pin_clk_14_, bottom_width_0_height_0_subtile_37__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__36_ccff_tail),
		.io_a2f_o(bottom_width_0_height_0_subtile_37__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_37__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__37_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__38 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[38]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[38]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[38]),
		.io_f2a_i(top_width_0_height_0_subtile_38__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_38__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_38__pin_clk_0_, bottom_width_0_height_0_subtile_38__pin_clk_1_, bottom_width_0_height_0_subtile_38__pin_clk_2_, bottom_width_0_height_0_subtile_38__pin_clk_3_, bottom_width_0_height_0_subtile_38__pin_clk_4_, bottom_width_0_height_0_subtile_38__pin_clk_5_, bottom_width_0_height_0_subtile_38__pin_clk_6_, bottom_width_0_height_0_subtile_38__pin_clk_7_, bottom_width_0_height_0_subtile_38__pin_clk_8_, bottom_width_0_height_0_subtile_38__pin_clk_9_, bottom_width_0_height_0_subtile_38__pin_clk_10_, bottom_width_0_height_0_subtile_38__pin_clk_11_, bottom_width_0_height_0_subtile_38__pin_clk_12_, bottom_width_0_height_0_subtile_38__pin_clk_13_, bottom_width_0_height_0_subtile_38__pin_clk_14_, bottom_width_0_height_0_subtile_38__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__37_ccff_tail),
		.io_a2f_o(bottom_width_0_height_0_subtile_38__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_38__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__38_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__39 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[39]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[39]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[39]),
		.io_f2a_i(top_width_0_height_0_subtile_39__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_39__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_39__pin_clk_0_, bottom_width_0_height_0_subtile_39__pin_clk_1_, bottom_width_0_height_0_subtile_39__pin_clk_2_, bottom_width_0_height_0_subtile_39__pin_clk_3_, bottom_width_0_height_0_subtile_39__pin_clk_4_, bottom_width_0_height_0_subtile_39__pin_clk_5_, bottom_width_0_height_0_subtile_39__pin_clk_6_, bottom_width_0_height_0_subtile_39__pin_clk_7_, bottom_width_0_height_0_subtile_39__pin_clk_8_, bottom_width_0_height_0_subtile_39__pin_clk_9_, bottom_width_0_height_0_subtile_39__pin_clk_10_, bottom_width_0_height_0_subtile_39__pin_clk_11_, bottom_width_0_height_0_subtile_39__pin_clk_12_, bottom_width_0_height_0_subtile_39__pin_clk_13_, bottom_width_0_height_0_subtile_39__pin_clk_14_, bottom_width_0_height_0_subtile_39__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__38_ccff_tail),
		.io_a2f_o(bottom_width_0_height_0_subtile_39__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_39__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__39_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__40 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[40]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[40]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[40]),
		.io_f2a_i(top_width_0_height_0_subtile_40__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_40__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_40__pin_clk_0_, bottom_width_0_height_0_subtile_40__pin_clk_1_, bottom_width_0_height_0_subtile_40__pin_clk_2_, bottom_width_0_height_0_subtile_40__pin_clk_3_, bottom_width_0_height_0_subtile_40__pin_clk_4_, bottom_width_0_height_0_subtile_40__pin_clk_5_, bottom_width_0_height_0_subtile_40__pin_clk_6_, bottom_width_0_height_0_subtile_40__pin_clk_7_, bottom_width_0_height_0_subtile_40__pin_clk_8_, bottom_width_0_height_0_subtile_40__pin_clk_9_, bottom_width_0_height_0_subtile_40__pin_clk_10_, bottom_width_0_height_0_subtile_40__pin_clk_11_, bottom_width_0_height_0_subtile_40__pin_clk_12_, bottom_width_0_height_0_subtile_40__pin_clk_13_, bottom_width_0_height_0_subtile_40__pin_clk_14_, bottom_width_0_height_0_subtile_40__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__39_ccff_tail),
		.io_a2f_o(bottom_width_0_height_0_subtile_40__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_40__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__40_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__41 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[41]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[41]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[41]),
		.io_f2a_i(top_width_0_height_0_subtile_41__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_41__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_41__pin_clk_0_, bottom_width_0_height_0_subtile_41__pin_clk_1_, bottom_width_0_height_0_subtile_41__pin_clk_2_, bottom_width_0_height_0_subtile_41__pin_clk_3_, bottom_width_0_height_0_subtile_41__pin_clk_4_, bottom_width_0_height_0_subtile_41__pin_clk_5_, bottom_width_0_height_0_subtile_41__pin_clk_6_, bottom_width_0_height_0_subtile_41__pin_clk_7_, bottom_width_0_height_0_subtile_41__pin_clk_8_, bottom_width_0_height_0_subtile_41__pin_clk_9_, bottom_width_0_height_0_subtile_41__pin_clk_10_, bottom_width_0_height_0_subtile_41__pin_clk_11_, bottom_width_0_height_0_subtile_41__pin_clk_12_, bottom_width_0_height_0_subtile_41__pin_clk_13_, bottom_width_0_height_0_subtile_41__pin_clk_14_, bottom_width_0_height_0_subtile_41__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__40_ccff_tail),
		.io_a2f_o(bottom_width_0_height_0_subtile_41__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_41__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__41_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__42 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[42]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[42]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[42]),
		.io_f2a_i(top_width_0_height_0_subtile_42__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_42__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_42__pin_clk_0_, bottom_width_0_height_0_subtile_42__pin_clk_1_, bottom_width_0_height_0_subtile_42__pin_clk_2_, bottom_width_0_height_0_subtile_42__pin_clk_3_, bottom_width_0_height_0_subtile_42__pin_clk_4_, bottom_width_0_height_0_subtile_42__pin_clk_5_, bottom_width_0_height_0_subtile_42__pin_clk_6_, bottom_width_0_height_0_subtile_42__pin_clk_7_, bottom_width_0_height_0_subtile_42__pin_clk_8_, bottom_width_0_height_0_subtile_42__pin_clk_9_, bottom_width_0_height_0_subtile_42__pin_clk_10_, bottom_width_0_height_0_subtile_42__pin_clk_11_, bottom_width_0_height_0_subtile_42__pin_clk_12_, bottom_width_0_height_0_subtile_42__pin_clk_13_, bottom_width_0_height_0_subtile_42__pin_clk_14_, bottom_width_0_height_0_subtile_42__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__41_ccff_tail),
		.io_a2f_o(bottom_width_0_height_0_subtile_42__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_42__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__42_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__43 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[43]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[43]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[43]),
		.io_f2a_i(top_width_0_height_0_subtile_43__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_43__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_43__pin_clk_0_, bottom_width_0_height_0_subtile_43__pin_clk_1_, bottom_width_0_height_0_subtile_43__pin_clk_2_, bottom_width_0_height_0_subtile_43__pin_clk_3_, bottom_width_0_height_0_subtile_43__pin_clk_4_, bottom_width_0_height_0_subtile_43__pin_clk_5_, bottom_width_0_height_0_subtile_43__pin_clk_6_, bottom_width_0_height_0_subtile_43__pin_clk_7_, bottom_width_0_height_0_subtile_43__pin_clk_8_, bottom_width_0_height_0_subtile_43__pin_clk_9_, bottom_width_0_height_0_subtile_43__pin_clk_10_, bottom_width_0_height_0_subtile_43__pin_clk_11_, bottom_width_0_height_0_subtile_43__pin_clk_12_, bottom_width_0_height_0_subtile_43__pin_clk_13_, bottom_width_0_height_0_subtile_43__pin_clk_14_, bottom_width_0_height_0_subtile_43__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__42_ccff_tail),
		.io_a2f_o(bottom_width_0_height_0_subtile_43__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_43__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__43_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__44 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[44]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[44]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[44]),
		.io_f2a_i(top_width_0_height_0_subtile_44__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_44__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_44__pin_clk_0_, bottom_width_0_height_0_subtile_44__pin_clk_1_, bottom_width_0_height_0_subtile_44__pin_clk_2_, bottom_width_0_height_0_subtile_44__pin_clk_3_, bottom_width_0_height_0_subtile_44__pin_clk_4_, bottom_width_0_height_0_subtile_44__pin_clk_5_, bottom_width_0_height_0_subtile_44__pin_clk_6_, bottom_width_0_height_0_subtile_44__pin_clk_7_, bottom_width_0_height_0_subtile_44__pin_clk_8_, bottom_width_0_height_0_subtile_44__pin_clk_9_, bottom_width_0_height_0_subtile_44__pin_clk_10_, bottom_width_0_height_0_subtile_44__pin_clk_11_, bottom_width_0_height_0_subtile_44__pin_clk_12_, bottom_width_0_height_0_subtile_44__pin_clk_13_, bottom_width_0_height_0_subtile_44__pin_clk_14_, bottom_width_0_height_0_subtile_44__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__43_ccff_tail),
		.io_a2f_o(bottom_width_0_height_0_subtile_44__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_44__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__44_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__45 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[45]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[45]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[45]),
		.io_f2a_i(top_width_0_height_0_subtile_45__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_45__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_45__pin_clk_0_, bottom_width_0_height_0_subtile_45__pin_clk_1_, bottom_width_0_height_0_subtile_45__pin_clk_2_, bottom_width_0_height_0_subtile_45__pin_clk_3_, bottom_width_0_height_0_subtile_45__pin_clk_4_, bottom_width_0_height_0_subtile_45__pin_clk_5_, bottom_width_0_height_0_subtile_45__pin_clk_6_, bottom_width_0_height_0_subtile_45__pin_clk_7_, bottom_width_0_height_0_subtile_45__pin_clk_8_, bottom_width_0_height_0_subtile_45__pin_clk_9_, bottom_width_0_height_0_subtile_45__pin_clk_10_, bottom_width_0_height_0_subtile_45__pin_clk_11_, bottom_width_0_height_0_subtile_45__pin_clk_12_, bottom_width_0_height_0_subtile_45__pin_clk_13_, bottom_width_0_height_0_subtile_45__pin_clk_14_, bottom_width_0_height_0_subtile_45__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__44_ccff_tail),
		.io_a2f_o(bottom_width_0_height_0_subtile_45__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_45__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__45_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__46 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[46]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[46]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[46]),
		.io_f2a_i(top_width_0_height_0_subtile_46__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_46__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_46__pin_clk_0_, bottom_width_0_height_0_subtile_46__pin_clk_1_, bottom_width_0_height_0_subtile_46__pin_clk_2_, bottom_width_0_height_0_subtile_46__pin_clk_3_, bottom_width_0_height_0_subtile_46__pin_clk_4_, bottom_width_0_height_0_subtile_46__pin_clk_5_, bottom_width_0_height_0_subtile_46__pin_clk_6_, bottom_width_0_height_0_subtile_46__pin_clk_7_, bottom_width_0_height_0_subtile_46__pin_clk_8_, bottom_width_0_height_0_subtile_46__pin_clk_9_, bottom_width_0_height_0_subtile_46__pin_clk_10_, bottom_width_0_height_0_subtile_46__pin_clk_11_, bottom_width_0_height_0_subtile_46__pin_clk_12_, bottom_width_0_height_0_subtile_46__pin_clk_13_, bottom_width_0_height_0_subtile_46__pin_clk_14_, bottom_width_0_height_0_subtile_46__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__45_ccff_tail),
		.io_a2f_o(bottom_width_0_height_0_subtile_46__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_46__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__46_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__47 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[47]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[47]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[47]),
		.io_f2a_i(top_width_0_height_0_subtile_47__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_47__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_47__pin_clk_0_, bottom_width_0_height_0_subtile_47__pin_clk_1_, bottom_width_0_height_0_subtile_47__pin_clk_2_, bottom_width_0_height_0_subtile_47__pin_clk_3_, bottom_width_0_height_0_subtile_47__pin_clk_4_, bottom_width_0_height_0_subtile_47__pin_clk_5_, bottom_width_0_height_0_subtile_47__pin_clk_6_, bottom_width_0_height_0_subtile_47__pin_clk_7_, bottom_width_0_height_0_subtile_47__pin_clk_8_, bottom_width_0_height_0_subtile_47__pin_clk_9_, bottom_width_0_height_0_subtile_47__pin_clk_10_, bottom_width_0_height_0_subtile_47__pin_clk_11_, bottom_width_0_height_0_subtile_47__pin_clk_12_, bottom_width_0_height_0_subtile_47__pin_clk_13_, bottom_width_0_height_0_subtile_47__pin_clk_14_, bottom_width_0_height_0_subtile_47__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__46_ccff_tail),
		.io_a2f_o(bottom_width_0_height_0_subtile_47__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_47__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__47_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__48 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[48]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[48]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[48]),
		.io_f2a_i(top_width_0_height_0_subtile_48__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_48__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_48__pin_clk_0_, bottom_width_0_height_0_subtile_48__pin_clk_1_, bottom_width_0_height_0_subtile_48__pin_clk_2_, bottom_width_0_height_0_subtile_48__pin_clk_3_, bottom_width_0_height_0_subtile_48__pin_clk_4_, bottom_width_0_height_0_subtile_48__pin_clk_5_, bottom_width_0_height_0_subtile_48__pin_clk_6_, bottom_width_0_height_0_subtile_48__pin_clk_7_, bottom_width_0_height_0_subtile_48__pin_clk_8_, bottom_width_0_height_0_subtile_48__pin_clk_9_, bottom_width_0_height_0_subtile_48__pin_clk_10_, bottom_width_0_height_0_subtile_48__pin_clk_11_, bottom_width_0_height_0_subtile_48__pin_clk_12_, bottom_width_0_height_0_subtile_48__pin_clk_13_, bottom_width_0_height_0_subtile_48__pin_clk_14_, bottom_width_0_height_0_subtile_48__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__47_ccff_tail),
		.io_a2f_o(bottom_width_0_height_0_subtile_48__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_48__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__48_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__49 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[49]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[49]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[49]),
		.io_f2a_i(top_width_0_height_0_subtile_49__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_49__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_49__pin_clk_0_, bottom_width_0_height_0_subtile_49__pin_clk_1_, bottom_width_0_height_0_subtile_49__pin_clk_2_, bottom_width_0_height_0_subtile_49__pin_clk_3_, bottom_width_0_height_0_subtile_49__pin_clk_4_, bottom_width_0_height_0_subtile_49__pin_clk_5_, bottom_width_0_height_0_subtile_49__pin_clk_6_, bottom_width_0_height_0_subtile_49__pin_clk_7_, bottom_width_0_height_0_subtile_49__pin_clk_8_, bottom_width_0_height_0_subtile_49__pin_clk_9_, bottom_width_0_height_0_subtile_49__pin_clk_10_, bottom_width_0_height_0_subtile_49__pin_clk_11_, bottom_width_0_height_0_subtile_49__pin_clk_12_, bottom_width_0_height_0_subtile_49__pin_clk_13_, bottom_width_0_height_0_subtile_49__pin_clk_14_, bottom_width_0_height_0_subtile_49__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__48_ccff_tail),
		.io_a2f_o(bottom_width_0_height_0_subtile_49__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_49__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__49_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__50 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[50]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[50]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[50]),
		.io_f2a_i(top_width_0_height_0_subtile_50__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_50__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_50__pin_clk_0_, bottom_width_0_height_0_subtile_50__pin_clk_1_, bottom_width_0_height_0_subtile_50__pin_clk_2_, bottom_width_0_height_0_subtile_50__pin_clk_3_, bottom_width_0_height_0_subtile_50__pin_clk_4_, bottom_width_0_height_0_subtile_50__pin_clk_5_, bottom_width_0_height_0_subtile_50__pin_clk_6_, bottom_width_0_height_0_subtile_50__pin_clk_7_, bottom_width_0_height_0_subtile_50__pin_clk_8_, bottom_width_0_height_0_subtile_50__pin_clk_9_, bottom_width_0_height_0_subtile_50__pin_clk_10_, bottom_width_0_height_0_subtile_50__pin_clk_11_, bottom_width_0_height_0_subtile_50__pin_clk_12_, bottom_width_0_height_0_subtile_50__pin_clk_13_, bottom_width_0_height_0_subtile_50__pin_clk_14_, bottom_width_0_height_0_subtile_50__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__49_ccff_tail),
		.io_a2f_o(bottom_width_0_height_0_subtile_50__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_50__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__50_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__51 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[51]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[51]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[51]),
		.io_f2a_i(top_width_0_height_0_subtile_51__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_51__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_51__pin_clk_0_, bottom_width_0_height_0_subtile_51__pin_clk_1_, bottom_width_0_height_0_subtile_51__pin_clk_2_, bottom_width_0_height_0_subtile_51__pin_clk_3_, bottom_width_0_height_0_subtile_51__pin_clk_4_, bottom_width_0_height_0_subtile_51__pin_clk_5_, bottom_width_0_height_0_subtile_51__pin_clk_6_, bottom_width_0_height_0_subtile_51__pin_clk_7_, bottom_width_0_height_0_subtile_51__pin_clk_8_, bottom_width_0_height_0_subtile_51__pin_clk_9_, bottom_width_0_height_0_subtile_51__pin_clk_10_, bottom_width_0_height_0_subtile_51__pin_clk_11_, bottom_width_0_height_0_subtile_51__pin_clk_12_, bottom_width_0_height_0_subtile_51__pin_clk_13_, bottom_width_0_height_0_subtile_51__pin_clk_14_, bottom_width_0_height_0_subtile_51__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__50_ccff_tail),
		.io_a2f_o(bottom_width_0_height_0_subtile_51__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_51__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__51_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__52 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[52]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[52]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[52]),
		.io_f2a_i(top_width_0_height_0_subtile_52__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_52__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_52__pin_clk_0_, bottom_width_0_height_0_subtile_52__pin_clk_1_, bottom_width_0_height_0_subtile_52__pin_clk_2_, bottom_width_0_height_0_subtile_52__pin_clk_3_, bottom_width_0_height_0_subtile_52__pin_clk_4_, bottom_width_0_height_0_subtile_52__pin_clk_5_, bottom_width_0_height_0_subtile_52__pin_clk_6_, bottom_width_0_height_0_subtile_52__pin_clk_7_, bottom_width_0_height_0_subtile_52__pin_clk_8_, bottom_width_0_height_0_subtile_52__pin_clk_9_, bottom_width_0_height_0_subtile_52__pin_clk_10_, bottom_width_0_height_0_subtile_52__pin_clk_11_, bottom_width_0_height_0_subtile_52__pin_clk_12_, bottom_width_0_height_0_subtile_52__pin_clk_13_, bottom_width_0_height_0_subtile_52__pin_clk_14_, bottom_width_0_height_0_subtile_52__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__51_ccff_tail),
		.io_a2f_o(bottom_width_0_height_0_subtile_52__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_52__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__52_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__53 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[53]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[53]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[53]),
		.io_f2a_i(top_width_0_height_0_subtile_53__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_53__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_53__pin_clk_0_, bottom_width_0_height_0_subtile_53__pin_clk_1_, bottom_width_0_height_0_subtile_53__pin_clk_2_, bottom_width_0_height_0_subtile_53__pin_clk_3_, bottom_width_0_height_0_subtile_53__pin_clk_4_, bottom_width_0_height_0_subtile_53__pin_clk_5_, bottom_width_0_height_0_subtile_53__pin_clk_6_, bottom_width_0_height_0_subtile_53__pin_clk_7_, bottom_width_0_height_0_subtile_53__pin_clk_8_, bottom_width_0_height_0_subtile_53__pin_clk_9_, bottom_width_0_height_0_subtile_53__pin_clk_10_, bottom_width_0_height_0_subtile_53__pin_clk_11_, bottom_width_0_height_0_subtile_53__pin_clk_12_, bottom_width_0_height_0_subtile_53__pin_clk_13_, bottom_width_0_height_0_subtile_53__pin_clk_14_, bottom_width_0_height_0_subtile_53__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__52_ccff_tail),
		.io_a2f_o(bottom_width_0_height_0_subtile_53__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_53__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__53_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__54 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[54]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[54]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[54]),
		.io_f2a_i(top_width_0_height_0_subtile_54__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_54__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_54__pin_clk_0_, bottom_width_0_height_0_subtile_54__pin_clk_1_, bottom_width_0_height_0_subtile_54__pin_clk_2_, bottom_width_0_height_0_subtile_54__pin_clk_3_, bottom_width_0_height_0_subtile_54__pin_clk_4_, bottom_width_0_height_0_subtile_54__pin_clk_5_, bottom_width_0_height_0_subtile_54__pin_clk_6_, bottom_width_0_height_0_subtile_54__pin_clk_7_, bottom_width_0_height_0_subtile_54__pin_clk_8_, bottom_width_0_height_0_subtile_54__pin_clk_9_, bottom_width_0_height_0_subtile_54__pin_clk_10_, bottom_width_0_height_0_subtile_54__pin_clk_11_, bottom_width_0_height_0_subtile_54__pin_clk_12_, bottom_width_0_height_0_subtile_54__pin_clk_13_, bottom_width_0_height_0_subtile_54__pin_clk_14_, bottom_width_0_height_0_subtile_54__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__53_ccff_tail),
		.io_a2f_o(bottom_width_0_height_0_subtile_54__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_54__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__54_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__55 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[55]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[55]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[55]),
		.io_f2a_i(top_width_0_height_0_subtile_55__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_55__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_55__pin_clk_0_, bottom_width_0_height_0_subtile_55__pin_clk_1_, bottom_width_0_height_0_subtile_55__pin_clk_2_, bottom_width_0_height_0_subtile_55__pin_clk_3_, bottom_width_0_height_0_subtile_55__pin_clk_4_, bottom_width_0_height_0_subtile_55__pin_clk_5_, bottom_width_0_height_0_subtile_55__pin_clk_6_, bottom_width_0_height_0_subtile_55__pin_clk_7_, bottom_width_0_height_0_subtile_55__pin_clk_8_, bottom_width_0_height_0_subtile_55__pin_clk_9_, bottom_width_0_height_0_subtile_55__pin_clk_10_, bottom_width_0_height_0_subtile_55__pin_clk_11_, bottom_width_0_height_0_subtile_55__pin_clk_12_, bottom_width_0_height_0_subtile_55__pin_clk_13_, bottom_width_0_height_0_subtile_55__pin_clk_14_, bottom_width_0_height_0_subtile_55__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__54_ccff_tail),
		.io_a2f_o(bottom_width_0_height_0_subtile_55__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_55__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__55_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__56 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[56]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[56]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[56]),
		.io_f2a_i(top_width_0_height_0_subtile_56__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_56__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_56__pin_clk_0_, bottom_width_0_height_0_subtile_56__pin_clk_1_, bottom_width_0_height_0_subtile_56__pin_clk_2_, bottom_width_0_height_0_subtile_56__pin_clk_3_, bottom_width_0_height_0_subtile_56__pin_clk_4_, bottom_width_0_height_0_subtile_56__pin_clk_5_, bottom_width_0_height_0_subtile_56__pin_clk_6_, bottom_width_0_height_0_subtile_56__pin_clk_7_, bottom_width_0_height_0_subtile_56__pin_clk_8_, bottom_width_0_height_0_subtile_56__pin_clk_9_, bottom_width_0_height_0_subtile_56__pin_clk_10_, bottom_width_0_height_0_subtile_56__pin_clk_11_, bottom_width_0_height_0_subtile_56__pin_clk_12_, bottom_width_0_height_0_subtile_56__pin_clk_13_, bottom_width_0_height_0_subtile_56__pin_clk_14_, bottom_width_0_height_0_subtile_56__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__55_ccff_tail),
		.io_a2f_o(bottom_width_0_height_0_subtile_56__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_56__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__56_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__57 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[57]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[57]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[57]),
		.io_f2a_i(top_width_0_height_0_subtile_57__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_57__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_57__pin_clk_0_, bottom_width_0_height_0_subtile_57__pin_clk_1_, bottom_width_0_height_0_subtile_57__pin_clk_2_, bottom_width_0_height_0_subtile_57__pin_clk_3_, bottom_width_0_height_0_subtile_57__pin_clk_4_, bottom_width_0_height_0_subtile_57__pin_clk_5_, bottom_width_0_height_0_subtile_57__pin_clk_6_, bottom_width_0_height_0_subtile_57__pin_clk_7_, bottom_width_0_height_0_subtile_57__pin_clk_8_, bottom_width_0_height_0_subtile_57__pin_clk_9_, bottom_width_0_height_0_subtile_57__pin_clk_10_, bottom_width_0_height_0_subtile_57__pin_clk_11_, bottom_width_0_height_0_subtile_57__pin_clk_12_, bottom_width_0_height_0_subtile_57__pin_clk_13_, bottom_width_0_height_0_subtile_57__pin_clk_14_, bottom_width_0_height_0_subtile_57__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__56_ccff_tail),
		.io_a2f_o(bottom_width_0_height_0_subtile_57__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_57__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__57_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__58 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[58]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[58]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[58]),
		.io_f2a_i(top_width_0_height_0_subtile_58__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_58__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_58__pin_clk_0_, bottom_width_0_height_0_subtile_58__pin_clk_1_, bottom_width_0_height_0_subtile_58__pin_clk_2_, bottom_width_0_height_0_subtile_58__pin_clk_3_, bottom_width_0_height_0_subtile_58__pin_clk_4_, bottom_width_0_height_0_subtile_58__pin_clk_5_, bottom_width_0_height_0_subtile_58__pin_clk_6_, bottom_width_0_height_0_subtile_58__pin_clk_7_, bottom_width_0_height_0_subtile_58__pin_clk_8_, bottom_width_0_height_0_subtile_58__pin_clk_9_, bottom_width_0_height_0_subtile_58__pin_clk_10_, bottom_width_0_height_0_subtile_58__pin_clk_11_, bottom_width_0_height_0_subtile_58__pin_clk_12_, bottom_width_0_height_0_subtile_58__pin_clk_13_, bottom_width_0_height_0_subtile_58__pin_clk_14_, bottom_width_0_height_0_subtile_58__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__57_ccff_tail),
		.io_a2f_o(bottom_width_0_height_0_subtile_58__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_58__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__58_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__59 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[59]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[59]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[59]),
		.io_f2a_i(top_width_0_height_0_subtile_59__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_59__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_59__pin_clk_0_, bottom_width_0_height_0_subtile_59__pin_clk_1_, bottom_width_0_height_0_subtile_59__pin_clk_2_, bottom_width_0_height_0_subtile_59__pin_clk_3_, bottom_width_0_height_0_subtile_59__pin_clk_4_, bottom_width_0_height_0_subtile_59__pin_clk_5_, bottom_width_0_height_0_subtile_59__pin_clk_6_, bottom_width_0_height_0_subtile_59__pin_clk_7_, bottom_width_0_height_0_subtile_59__pin_clk_8_, bottom_width_0_height_0_subtile_59__pin_clk_9_, bottom_width_0_height_0_subtile_59__pin_clk_10_, bottom_width_0_height_0_subtile_59__pin_clk_11_, bottom_width_0_height_0_subtile_59__pin_clk_12_, bottom_width_0_height_0_subtile_59__pin_clk_13_, bottom_width_0_height_0_subtile_59__pin_clk_14_, bottom_width_0_height_0_subtile_59__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__58_ccff_tail),
		.io_a2f_o(bottom_width_0_height_0_subtile_59__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_59__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__59_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__60 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[60]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[60]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[60]),
		.io_f2a_i(top_width_0_height_0_subtile_60__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_60__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_60__pin_clk_0_, bottom_width_0_height_0_subtile_60__pin_clk_1_, bottom_width_0_height_0_subtile_60__pin_clk_2_, bottom_width_0_height_0_subtile_60__pin_clk_3_, bottom_width_0_height_0_subtile_60__pin_clk_4_, bottom_width_0_height_0_subtile_60__pin_clk_5_, bottom_width_0_height_0_subtile_60__pin_clk_6_, bottom_width_0_height_0_subtile_60__pin_clk_7_, bottom_width_0_height_0_subtile_60__pin_clk_8_, bottom_width_0_height_0_subtile_60__pin_clk_9_, bottom_width_0_height_0_subtile_60__pin_clk_10_, bottom_width_0_height_0_subtile_60__pin_clk_11_, bottom_width_0_height_0_subtile_60__pin_clk_12_, bottom_width_0_height_0_subtile_60__pin_clk_13_, bottom_width_0_height_0_subtile_60__pin_clk_14_, bottom_width_0_height_0_subtile_60__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__59_ccff_tail),
		.io_a2f_o(bottom_width_0_height_0_subtile_60__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_60__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__60_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__61 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[61]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[61]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[61]),
		.io_f2a_i(top_width_0_height_0_subtile_61__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_61__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_61__pin_clk_0_, bottom_width_0_height_0_subtile_61__pin_clk_1_, bottom_width_0_height_0_subtile_61__pin_clk_2_, bottom_width_0_height_0_subtile_61__pin_clk_3_, bottom_width_0_height_0_subtile_61__pin_clk_4_, bottom_width_0_height_0_subtile_61__pin_clk_5_, bottom_width_0_height_0_subtile_61__pin_clk_6_, bottom_width_0_height_0_subtile_61__pin_clk_7_, bottom_width_0_height_0_subtile_61__pin_clk_8_, bottom_width_0_height_0_subtile_61__pin_clk_9_, bottom_width_0_height_0_subtile_61__pin_clk_10_, bottom_width_0_height_0_subtile_61__pin_clk_11_, bottom_width_0_height_0_subtile_61__pin_clk_12_, bottom_width_0_height_0_subtile_61__pin_clk_13_, bottom_width_0_height_0_subtile_61__pin_clk_14_, bottom_width_0_height_0_subtile_61__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__60_ccff_tail),
		.io_a2f_o(bottom_width_0_height_0_subtile_61__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_61__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__61_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__62 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[62]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[62]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[62]),
		.io_f2a_i(top_width_0_height_0_subtile_62__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_62__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_62__pin_clk_0_, bottom_width_0_height_0_subtile_62__pin_clk_1_, bottom_width_0_height_0_subtile_62__pin_clk_2_, bottom_width_0_height_0_subtile_62__pin_clk_3_, bottom_width_0_height_0_subtile_62__pin_clk_4_, bottom_width_0_height_0_subtile_62__pin_clk_5_, bottom_width_0_height_0_subtile_62__pin_clk_6_, bottom_width_0_height_0_subtile_62__pin_clk_7_, bottom_width_0_height_0_subtile_62__pin_clk_8_, bottom_width_0_height_0_subtile_62__pin_clk_9_, bottom_width_0_height_0_subtile_62__pin_clk_10_, bottom_width_0_height_0_subtile_62__pin_clk_11_, bottom_width_0_height_0_subtile_62__pin_clk_12_, bottom_width_0_height_0_subtile_62__pin_clk_13_, bottom_width_0_height_0_subtile_62__pin_clk_14_, bottom_width_0_height_0_subtile_62__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__61_ccff_tail),
		.io_a2f_o(bottom_width_0_height_0_subtile_62__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_62__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__62_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__63 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[63]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[63]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[63]),
		.io_f2a_i(top_width_0_height_0_subtile_63__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_63__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_63__pin_clk_0_, bottom_width_0_height_0_subtile_63__pin_clk_1_, bottom_width_0_height_0_subtile_63__pin_clk_2_, bottom_width_0_height_0_subtile_63__pin_clk_3_, bottom_width_0_height_0_subtile_63__pin_clk_4_, bottom_width_0_height_0_subtile_63__pin_clk_5_, bottom_width_0_height_0_subtile_63__pin_clk_6_, bottom_width_0_height_0_subtile_63__pin_clk_7_, bottom_width_0_height_0_subtile_63__pin_clk_8_, bottom_width_0_height_0_subtile_63__pin_clk_9_, bottom_width_0_height_0_subtile_63__pin_clk_10_, bottom_width_0_height_0_subtile_63__pin_clk_11_, bottom_width_0_height_0_subtile_63__pin_clk_12_, bottom_width_0_height_0_subtile_63__pin_clk_13_, bottom_width_0_height_0_subtile_63__pin_clk_14_, bottom_width_0_height_0_subtile_63__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__62_ccff_tail),
		.io_a2f_o(bottom_width_0_height_0_subtile_63__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_63__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__63_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__64 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[64]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[64]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[64]),
		.io_f2a_i(top_width_0_height_0_subtile_64__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_64__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_64__pin_clk_0_, bottom_width_0_height_0_subtile_64__pin_clk_1_, bottom_width_0_height_0_subtile_64__pin_clk_2_, bottom_width_0_height_0_subtile_64__pin_clk_3_, bottom_width_0_height_0_subtile_64__pin_clk_4_, bottom_width_0_height_0_subtile_64__pin_clk_5_, bottom_width_0_height_0_subtile_64__pin_clk_6_, bottom_width_0_height_0_subtile_64__pin_clk_7_, bottom_width_0_height_0_subtile_64__pin_clk_8_, bottom_width_0_height_0_subtile_64__pin_clk_9_, bottom_width_0_height_0_subtile_64__pin_clk_10_, bottom_width_0_height_0_subtile_64__pin_clk_11_, bottom_width_0_height_0_subtile_64__pin_clk_12_, bottom_width_0_height_0_subtile_64__pin_clk_13_, bottom_width_0_height_0_subtile_64__pin_clk_14_, bottom_width_0_height_0_subtile_64__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__63_ccff_tail),
		.io_a2f_o(bottom_width_0_height_0_subtile_64__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_64__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__64_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__65 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[65]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[65]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[65]),
		.io_f2a_i(top_width_0_height_0_subtile_65__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_65__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_65__pin_clk_0_, bottom_width_0_height_0_subtile_65__pin_clk_1_, bottom_width_0_height_0_subtile_65__pin_clk_2_, bottom_width_0_height_0_subtile_65__pin_clk_3_, bottom_width_0_height_0_subtile_65__pin_clk_4_, bottom_width_0_height_0_subtile_65__pin_clk_5_, bottom_width_0_height_0_subtile_65__pin_clk_6_, bottom_width_0_height_0_subtile_65__pin_clk_7_, bottom_width_0_height_0_subtile_65__pin_clk_8_, bottom_width_0_height_0_subtile_65__pin_clk_9_, bottom_width_0_height_0_subtile_65__pin_clk_10_, bottom_width_0_height_0_subtile_65__pin_clk_11_, bottom_width_0_height_0_subtile_65__pin_clk_12_, bottom_width_0_height_0_subtile_65__pin_clk_13_, bottom_width_0_height_0_subtile_65__pin_clk_14_, bottom_width_0_height_0_subtile_65__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__64_ccff_tail),
		.io_a2f_o(bottom_width_0_height_0_subtile_65__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_65__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__65_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__66 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[66]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[66]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[66]),
		.io_f2a_i(top_width_0_height_0_subtile_66__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_66__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_66__pin_clk_0_, bottom_width_0_height_0_subtile_66__pin_clk_1_, bottom_width_0_height_0_subtile_66__pin_clk_2_, bottom_width_0_height_0_subtile_66__pin_clk_3_, bottom_width_0_height_0_subtile_66__pin_clk_4_, bottom_width_0_height_0_subtile_66__pin_clk_5_, bottom_width_0_height_0_subtile_66__pin_clk_6_, bottom_width_0_height_0_subtile_66__pin_clk_7_, bottom_width_0_height_0_subtile_66__pin_clk_8_, bottom_width_0_height_0_subtile_66__pin_clk_9_, bottom_width_0_height_0_subtile_66__pin_clk_10_, bottom_width_0_height_0_subtile_66__pin_clk_11_, bottom_width_0_height_0_subtile_66__pin_clk_12_, bottom_width_0_height_0_subtile_66__pin_clk_13_, bottom_width_0_height_0_subtile_66__pin_clk_14_, bottom_width_0_height_0_subtile_66__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__65_ccff_tail),
		.io_a2f_o(bottom_width_0_height_0_subtile_66__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_66__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__66_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__67 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[67]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[67]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[67]),
		.io_f2a_i(top_width_0_height_0_subtile_67__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_67__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_67__pin_clk_0_, bottom_width_0_height_0_subtile_67__pin_clk_1_, bottom_width_0_height_0_subtile_67__pin_clk_2_, bottom_width_0_height_0_subtile_67__pin_clk_3_, bottom_width_0_height_0_subtile_67__pin_clk_4_, bottom_width_0_height_0_subtile_67__pin_clk_5_, bottom_width_0_height_0_subtile_67__pin_clk_6_, bottom_width_0_height_0_subtile_67__pin_clk_7_, bottom_width_0_height_0_subtile_67__pin_clk_8_, bottom_width_0_height_0_subtile_67__pin_clk_9_, bottom_width_0_height_0_subtile_67__pin_clk_10_, bottom_width_0_height_0_subtile_67__pin_clk_11_, bottom_width_0_height_0_subtile_67__pin_clk_12_, bottom_width_0_height_0_subtile_67__pin_clk_13_, bottom_width_0_height_0_subtile_67__pin_clk_14_, bottom_width_0_height_0_subtile_67__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__66_ccff_tail),
		.io_a2f_o(bottom_width_0_height_0_subtile_67__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_67__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__67_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__68 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[68]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[68]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[68]),
		.io_f2a_i(top_width_0_height_0_subtile_68__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_68__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_68__pin_clk_0_, bottom_width_0_height_0_subtile_68__pin_clk_1_, bottom_width_0_height_0_subtile_68__pin_clk_2_, bottom_width_0_height_0_subtile_68__pin_clk_3_, bottom_width_0_height_0_subtile_68__pin_clk_4_, bottom_width_0_height_0_subtile_68__pin_clk_5_, bottom_width_0_height_0_subtile_68__pin_clk_6_, bottom_width_0_height_0_subtile_68__pin_clk_7_, bottom_width_0_height_0_subtile_68__pin_clk_8_, bottom_width_0_height_0_subtile_68__pin_clk_9_, bottom_width_0_height_0_subtile_68__pin_clk_10_, bottom_width_0_height_0_subtile_68__pin_clk_11_, bottom_width_0_height_0_subtile_68__pin_clk_12_, bottom_width_0_height_0_subtile_68__pin_clk_13_, bottom_width_0_height_0_subtile_68__pin_clk_14_, bottom_width_0_height_0_subtile_68__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__67_ccff_tail),
		.io_a2f_o(bottom_width_0_height_0_subtile_68__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_68__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__68_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__69 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[69]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[69]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[69]),
		.io_f2a_i(top_width_0_height_0_subtile_69__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_69__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_69__pin_clk_0_, bottom_width_0_height_0_subtile_69__pin_clk_1_, bottom_width_0_height_0_subtile_69__pin_clk_2_, bottom_width_0_height_0_subtile_69__pin_clk_3_, bottom_width_0_height_0_subtile_69__pin_clk_4_, bottom_width_0_height_0_subtile_69__pin_clk_5_, bottom_width_0_height_0_subtile_69__pin_clk_6_, bottom_width_0_height_0_subtile_69__pin_clk_7_, bottom_width_0_height_0_subtile_69__pin_clk_8_, bottom_width_0_height_0_subtile_69__pin_clk_9_, bottom_width_0_height_0_subtile_69__pin_clk_10_, bottom_width_0_height_0_subtile_69__pin_clk_11_, bottom_width_0_height_0_subtile_69__pin_clk_12_, bottom_width_0_height_0_subtile_69__pin_clk_13_, bottom_width_0_height_0_subtile_69__pin_clk_14_, bottom_width_0_height_0_subtile_69__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__68_ccff_tail),
		.io_a2f_o(bottom_width_0_height_0_subtile_69__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_69__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__69_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__70 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[70]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[70]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[70]),
		.io_f2a_i(top_width_0_height_0_subtile_70__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_70__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_70__pin_clk_0_, bottom_width_0_height_0_subtile_70__pin_clk_1_, bottom_width_0_height_0_subtile_70__pin_clk_2_, bottom_width_0_height_0_subtile_70__pin_clk_3_, bottom_width_0_height_0_subtile_70__pin_clk_4_, bottom_width_0_height_0_subtile_70__pin_clk_5_, bottom_width_0_height_0_subtile_70__pin_clk_6_, bottom_width_0_height_0_subtile_70__pin_clk_7_, bottom_width_0_height_0_subtile_70__pin_clk_8_, bottom_width_0_height_0_subtile_70__pin_clk_9_, bottom_width_0_height_0_subtile_70__pin_clk_10_, bottom_width_0_height_0_subtile_70__pin_clk_11_, bottom_width_0_height_0_subtile_70__pin_clk_12_, bottom_width_0_height_0_subtile_70__pin_clk_13_, bottom_width_0_height_0_subtile_70__pin_clk_14_, bottom_width_0_height_0_subtile_70__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__69_ccff_tail),
		.io_a2f_o(bottom_width_0_height_0_subtile_70__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_70__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_mode_io__70_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__71 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[71]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[71]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[71]),
		.io_f2a_i(top_width_0_height_0_subtile_71__pin_f2a_i_0_),
		.io_sc_in(left_width_0_height_0_subtile_71__pin_sc_in_0_),
		.io_clk({bottom_width_0_height_0_subtile_71__pin_clk_0_, bottom_width_0_height_0_subtile_71__pin_clk_1_, bottom_width_0_height_0_subtile_71__pin_clk_2_, bottom_width_0_height_0_subtile_71__pin_clk_3_, bottom_width_0_height_0_subtile_71__pin_clk_4_, bottom_width_0_height_0_subtile_71__pin_clk_5_, bottom_width_0_height_0_subtile_71__pin_clk_6_, bottom_width_0_height_0_subtile_71__pin_clk_7_, bottom_width_0_height_0_subtile_71__pin_clk_8_, bottom_width_0_height_0_subtile_71__pin_clk_9_, bottom_width_0_height_0_subtile_71__pin_clk_10_, bottom_width_0_height_0_subtile_71__pin_clk_11_, bottom_width_0_height_0_subtile_71__pin_clk_12_, bottom_width_0_height_0_subtile_71__pin_clk_13_, bottom_width_0_height_0_subtile_71__pin_clk_14_, bottom_width_0_height_0_subtile_71__pin_clk_15_}),
		.ccff_head(logical_tile_io_mode_io__70_ccff_tail),
		.io_a2f_o(bottom_width_0_height_0_subtile_71__pin_a2f_o_0_),
		.io_sc_out(left_width_0_height_0_subtile_71__pin_sc_out_0_),
		.ccff_tail(ccff_tail));

endmodule
// ----- END Verilog module for grid_io_bottom -----

//----- Default net type -----
`default_nettype none



// ----- END Grid Verilog module: grid_io_bottom -----

