module MultiplierLUT(a, b, z);
    input [1:0] a;
    input [1:0] b;
    output reg [3:0] z;

    always @(a, b) begin
        case ({a, b})
            4'b0000: z <= 4'b0000; // 0 * 0 = 0
            4'b0001: z <= 4'b0000; // 0 * 1 = 0
            4'b0010: z <= 4'b0000; // 0 * 2 = 0
            4'b0011: z <= 4'b0000; // 0 * 3 = 0
            4'b0100: z <= 4'b0000; // 1 * 0 = 0
            4'b0101: z <= 4'b0001; // 1 * 1 = 1
            4'b0110: z <= 4'b0010; // 1 * 2 = 2
            4'b0111: z <= 4'b0011; // 1 * 3 = 3
            4'b1000: z <= 4'b0000; // 2 * 0 = 0
            4'b1001: z <= 4'b0010; // 2 * 1 = 2
            4'b1010: z <= 4'b0100; // 2 * 2 = 4
            4'b1011: z <= 4'b0110; // 2 * 3 = 6
            4'b1100: z <= 4'b0000; // 3 * 0 = 0
            4'b1101: z <= 4'b0011; // 3 * 1 = 3
            4'b1110: z <= 4'b0110; // 3 * 2 = 6
            4'b1111: z <= 4'b1001; // 3 * 3 = 9
            default: z <= 0;
        endcase
    end
endmodule
