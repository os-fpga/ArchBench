//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for Unique Switch Blocks[2][0]
//	Author: Xifan TANG
//	Organization: University of Utah
//-------------------------------------------
//----- Time scale -----
`timescale 1ns / 1ps

//----- Default net type -----
`default_nettype wire

// ----- Verilog module for sb_2__0_ -----
module sb_2__0_(config_enable,
                prog_clock,
                chany_top_in,
                chanx_right_in,
                chanx_left_in,
                ccff_head,
                chany_top_out,
                chanx_right_out,
                chanx_left_out,
                ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_clock;
//----- INPUT PORTS -----
input [0:95] chany_top_in;
//----- INPUT PORTS -----
input [0:95] chanx_right_in;
//----- INPUT PORTS -----
input [0:95] chanx_left_in;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:95] chany_top_out;
//----- OUTPUT PORTS -----
output [0:95] chanx_right_out;
//----- OUTPUT PORTS -----
output [0:95] chanx_left_out;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:1] mux_tree_tapbuf_L1SB_size3_0_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size3_0_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size3_10_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size3_10_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size3_11_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size3_11_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size3_12_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size3_12_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size3_13_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size3_13_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size3_14_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size3_14_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size3_15_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size3_15_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size3_16_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size3_16_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size3_17_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size3_17_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size3_18_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size3_18_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size3_1_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size3_1_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size3_2_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size3_2_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size3_3_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size3_3_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size3_4_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size3_4_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size3_5_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size3_5_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size3_6_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size3_6_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size3_7_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size3_7_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size3_8_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size3_8_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size3_9_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size3_9_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_0_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_0_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_10_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_10_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_11_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_11_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_12_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_12_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_13_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_13_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_14_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_14_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_15_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_15_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_16_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_16_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_17_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_17_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_18_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_18_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_19_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_19_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_1_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_1_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_2_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_2_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_3_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_3_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_4_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_4_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_5_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_5_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_6_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_6_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_7_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_7_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_8_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_8_sram_inv;
wire [0:1] mux_tree_tapbuf_L1SB_size4_9_sram;
wire [0:1] mux_tree_tapbuf_L1SB_size4_9_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size5_0_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size5_0_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size5_10_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size5_10_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size5_11_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size5_11_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size5_12_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size5_12_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size5_13_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size5_13_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size5_14_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size5_14_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size5_15_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size5_15_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size5_16_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size5_16_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size5_17_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size5_17_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size5_1_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size5_1_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size5_2_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size5_2_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size5_3_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size5_3_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size5_4_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size5_4_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size5_5_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size5_5_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size5_6_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size5_6_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size5_7_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size5_7_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size5_8_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size5_8_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size5_9_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size5_9_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_0_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_0_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_10_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_10_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_11_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_11_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_12_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_12_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_13_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_13_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_14_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_14_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_15_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_15_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_16_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_16_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_17_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_17_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_18_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_18_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_19_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_19_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_1_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_1_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_20_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_20_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_21_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_21_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_22_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_22_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_23_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_23_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_24_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_24_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_25_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_25_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_26_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_26_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_27_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_27_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_28_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_28_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_29_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_29_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_2_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_2_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_30_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_30_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_31_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_31_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_32_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_32_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_33_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_33_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_34_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_34_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_35_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_35_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_36_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_36_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_37_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_37_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_38_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_38_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_39_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_39_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_3_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_3_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_40_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_40_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_41_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_41_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_4_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_4_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_5_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_5_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_6_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_6_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_7_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_7_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_8_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_8_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_9_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_9_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_0_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_0_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_10_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_10_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_11_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_11_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_12_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_12_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_13_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_13_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_14_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_14_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_15_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_15_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_16_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_16_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_1_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_1_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_2_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_2_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_3_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_3_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_4_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_4_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_5_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_5_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_6_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_6_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_7_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_7_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_8_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_8_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size4_9_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size4_9_sram_inv;

// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 115 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[20] = chanx_right_in[19];
// ----- Local connection due to Wire 116 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[21] = chanx_right_in[20];
// ----- Local connection due to Wire 117 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[22] = chanx_right_in[21];
// ----- Local connection due to Wire 119 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[24] = chanx_right_in[23];
// ----- Local connection due to Wire 120 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[25] = chanx_right_in[24];
// ----- Local connection due to Wire 121 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[26] = chanx_right_in[25];
// ----- Local connection due to Wire 123 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[28] = chanx_right_in[27];
// ----- Local connection due to Wire 124 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[29] = chanx_right_in[28];
// ----- Local connection due to Wire 125 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[30] = chanx_right_in[29];
// ----- Local connection due to Wire 127 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[32] = chanx_right_in[31];
// ----- Local connection due to Wire 128 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[33] = chanx_right_in[32];
// ----- Local connection due to Wire 129 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[34] = chanx_right_in[33];
// ----- Local connection due to Wire 131 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[36] = chanx_right_in[35];
// ----- Local connection due to Wire 132 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[37] = chanx_right_in[36];
// ----- Local connection due to Wire 133 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[38] = chanx_right_in[37];
// ----- Local connection due to Wire 135 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[40] = chanx_right_in[39];
// ----- Local connection due to Wire 136 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[41] = chanx_right_in[40];
// ----- Local connection due to Wire 137 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[42] = chanx_right_in[41];
// ----- Local connection due to Wire 139 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[44] = chanx_right_in[43];
// ----- Local connection due to Wire 140 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[45] = chanx_right_in[44];
// ----- Local connection due to Wire 141 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[46] = chanx_right_in[45];
// ----- Local connection due to Wire 143 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[48] = chanx_right_in[47];
// ----- Local connection due to Wire 144 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[49] = chanx_right_in[48];
// ----- Local connection due to Wire 145 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[50] = chanx_right_in[49];
// ----- Local connection due to Wire 147 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[52] = chanx_right_in[51];
// ----- Local connection due to Wire 148 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[53] = chanx_right_in[52];
// ----- Local connection due to Wire 149 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[54] = chanx_right_in[53];
// ----- Local connection due to Wire 151 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[56] = chanx_right_in[55];
// ----- Local connection due to Wire 152 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[57] = chanx_right_in[56];
// ----- Local connection due to Wire 153 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[58] = chanx_right_in[57];
// ----- Local connection due to Wire 155 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[60] = chanx_right_in[59];
// ----- Local connection due to Wire 156 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[61] = chanx_right_in[60];
// ----- Local connection due to Wire 157 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[62] = chanx_right_in[61];
// ----- Local connection due to Wire 159 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[64] = chanx_right_in[63];
// ----- Local connection due to Wire 160 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[65] = chanx_right_in[64];
// ----- Local connection due to Wire 161 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[66] = chanx_right_in[65];
// ----- Local connection due to Wire 163 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[68] = chanx_right_in[67];
// ----- Local connection due to Wire 164 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[69] = chanx_right_in[68];
// ----- Local connection due to Wire 165 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[70] = chanx_right_in[69];
// ----- Local connection due to Wire 167 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[72] = chanx_right_in[71];
// ----- Local connection due to Wire 168 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[73] = chanx_right_in[72];
// ----- Local connection due to Wire 169 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[74] = chanx_right_in[73];
// ----- Local connection due to Wire 171 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[76] = chanx_right_in[75];
// ----- Local connection due to Wire 172 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[77] = chanx_right_in[76];
// ----- Local connection due to Wire 173 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[78] = chanx_right_in[77];
// ----- Local connection due to Wire 175 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[80] = chanx_right_in[79];
// ----- Local connection due to Wire 176 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[81] = chanx_right_in[80];
// ----- Local connection due to Wire 177 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[82] = chanx_right_in[81];
// ----- Local connection due to Wire 179 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[84] = chanx_right_in[83];
// ----- Local connection due to Wire 180 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[85] = chanx_right_in[84];
// ----- Local connection due to Wire 181 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[86] = chanx_right_in[85];
// ----- Local connection due to Wire 183 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[88] = chanx_right_in[87];
// ----- Local connection due to Wire 184 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[89] = chanx_right_in[88];
// ----- Local connection due to Wire 185 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[90] = chanx_right_in[89];
// ----- Local connection due to Wire 187 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[92] = chanx_right_in[91];
// ----- Local connection due to Wire 188 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[93] = chanx_right_in[92];
// ----- Local connection due to Wire 189 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[94] = chanx_right_in[93];
// ----- Local connection due to Wire 194 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[94] = chanx_left_in[2];
// ----- Local connection due to Wire 195 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[93] = chanx_left_in[3];
// ----- Local connection due to Wire 196 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[92] = chanx_left_in[4];
// ----- Local connection due to Wire 197 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[91] = chanx_left_in[5];
// ----- Local connection due to Wire 198 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[90] = chanx_left_in[6];
// ----- Local connection due to Wire 199 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[89] = chanx_left_in[7];
// ----- Local connection due to Wire 200 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[88] = chanx_left_in[8];
// ----- Local connection due to Wire 201 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[87] = chanx_left_in[9];
// ----- Local connection due to Wire 202 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[86] = chanx_left_in[10];
// ----- Local connection due to Wire 203 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[85] = chanx_left_in[11];
// ----- Local connection due to Wire 204 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[84] = chanx_left_in[12];
// ----- Local connection due to Wire 205 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[83] = chanx_left_in[13];
// ----- Local connection due to Wire 206 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[82] = chanx_left_in[14];
// ----- Local connection due to Wire 207 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[81] = chanx_left_in[15];
// ----- Local connection due to Wire 208 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[80] = chanx_left_in[16];
// ----- Local connection due to Wire 209 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[79] = chanx_left_in[17];
// ----- Local connection due to Wire 210 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[78] = chanx_left_in[18];
// ----- Local connection due to Wire 211 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[20] = chanx_left_in[19];
// ----- Local connection due to Wire 212 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[21] = chanx_left_in[20];
// ----- Local connection due to Wire 213 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[22] = chanx_left_in[21];
// ----- Local connection due to Wire 214 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[77] = chanx_left_in[22];
// ----- Local connection due to Wire 215 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[24] = chanx_left_in[23];
// ----- Local connection due to Wire 216 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[25] = chanx_left_in[24];
// ----- Local connection due to Wire 217 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[26] = chanx_left_in[25];
// ----- Local connection due to Wire 218 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[76] = chanx_left_in[26];
// ----- Local connection due to Wire 219 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[28] = chanx_left_in[27];
// ----- Local connection due to Wire 220 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[29] = chanx_left_in[28];
// ----- Local connection due to Wire 221 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[30] = chanx_left_in[29];
// ----- Local connection due to Wire 222 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[75] = chanx_left_in[30];
// ----- Local connection due to Wire 223 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[32] = chanx_left_in[31];
// ----- Local connection due to Wire 224 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[33] = chanx_left_in[32];
// ----- Local connection due to Wire 225 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[34] = chanx_left_in[33];
// ----- Local connection due to Wire 226 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[74] = chanx_left_in[34];
// ----- Local connection due to Wire 227 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[36] = chanx_left_in[35];
// ----- Local connection due to Wire 228 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[37] = chanx_left_in[36];
// ----- Local connection due to Wire 229 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[38] = chanx_left_in[37];
// ----- Local connection due to Wire 230 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[73] = chanx_left_in[38];
// ----- Local connection due to Wire 231 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[40] = chanx_left_in[39];
// ----- Local connection due to Wire 232 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[41] = chanx_left_in[40];
// ----- Local connection due to Wire 233 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[42] = chanx_left_in[41];
// ----- Local connection due to Wire 234 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[72] = chanx_left_in[42];
// ----- Local connection due to Wire 235 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[44] = chanx_left_in[43];
// ----- Local connection due to Wire 236 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[45] = chanx_left_in[44];
// ----- Local connection due to Wire 237 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[46] = chanx_left_in[45];
// ----- Local connection due to Wire 238 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[71] = chanx_left_in[46];
// ----- Local connection due to Wire 239 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[48] = chanx_left_in[47];
// ----- Local connection due to Wire 240 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[49] = chanx_left_in[48];
// ----- Local connection due to Wire 241 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[50] = chanx_left_in[49];
// ----- Local connection due to Wire 242 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[70] = chanx_left_in[50];
// ----- Local connection due to Wire 243 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[52] = chanx_left_in[51];
// ----- Local connection due to Wire 244 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[53] = chanx_left_in[52];
// ----- Local connection due to Wire 245 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[54] = chanx_left_in[53];
// ----- Local connection due to Wire 246 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[69] = chanx_left_in[54];
// ----- Local connection due to Wire 247 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[56] = chanx_left_in[55];
// ----- Local connection due to Wire 248 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[57] = chanx_left_in[56];
// ----- Local connection due to Wire 249 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[58] = chanx_left_in[57];
// ----- Local connection due to Wire 250 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[68] = chanx_left_in[58];
// ----- Local connection due to Wire 251 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[60] = chanx_left_in[59];
// ----- Local connection due to Wire 252 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[61] = chanx_left_in[60];
// ----- Local connection due to Wire 253 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[62] = chanx_left_in[61];
// ----- Local connection due to Wire 254 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[67] = chanx_left_in[62];
// ----- Local connection due to Wire 255 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[64] = chanx_left_in[63];
// ----- Local connection due to Wire 256 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[65] = chanx_left_in[64];
// ----- Local connection due to Wire 257 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[66] = chanx_left_in[65];
// ----- Local connection due to Wire 258 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[66] = chanx_left_in[66];
// ----- Local connection due to Wire 259 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[68] = chanx_left_in[67];
// ----- Local connection due to Wire 260 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[69] = chanx_left_in[68];
// ----- Local connection due to Wire 261 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[70] = chanx_left_in[69];
// ----- Local connection due to Wire 262 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[65] = chanx_left_in[70];
// ----- Local connection due to Wire 263 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[72] = chanx_left_in[71];
// ----- Local connection due to Wire 264 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[73] = chanx_left_in[72];
// ----- Local connection due to Wire 265 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[74] = chanx_left_in[73];
// ----- Local connection due to Wire 266 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[64] = chanx_left_in[74];
// ----- Local connection due to Wire 267 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[76] = chanx_left_in[75];
// ----- Local connection due to Wire 268 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[77] = chanx_left_in[76];
// ----- Local connection due to Wire 269 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[78] = chanx_left_in[77];
// ----- Local connection due to Wire 270 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[63] = chanx_left_in[78];
// ----- Local connection due to Wire 271 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[80] = chanx_left_in[79];
// ----- Local connection due to Wire 272 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[81] = chanx_left_in[80];
// ----- Local connection due to Wire 273 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[82] = chanx_left_in[81];
// ----- Local connection due to Wire 274 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[62] = chanx_left_in[82];
// ----- Local connection due to Wire 275 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[84] = chanx_left_in[83];
// ----- Local connection due to Wire 276 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[85] = chanx_left_in[84];
// ----- Local connection due to Wire 277 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[86] = chanx_left_in[85];
// ----- Local connection due to Wire 278 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[61] = chanx_left_in[86];
// ----- Local connection due to Wire 279 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[88] = chanx_left_in[87];
// ----- Local connection due to Wire 280 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[89] = chanx_left_in[88];
// ----- Local connection due to Wire 281 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[90] = chanx_left_in[89];
// ----- Local connection due to Wire 282 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[60] = chanx_left_in[90];
// ----- Local connection due to Wire 283 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[92] = chanx_left_in[91];
// ----- Local connection due to Wire 284 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[93] = chanx_left_in[92];
// ----- Local connection due to Wire 285 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[94] = chanx_left_in[93];
// ----- Local connection due to Wire 286 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[59] = chanx_left_in[94];
// ----- Local connection due to Wire 287 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[58] = chanx_left_in[95];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	mux_tree_tapbuf_L1SB_size4 mux_top_track_0 (
		.in({chanx_right_in[1], chanx_right_in[19], chanx_left_in[0], chanx_left_in[19]}),
		.sram(mux_tree_tapbuf_L1SB_size4_0_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_0_sram_inv[0:1]),
		.out(chany_top_out[0]));

	mux_tree_tapbuf_L1SB_size4 mux_right_track_0 (
		.in({chany_top_in[38], chany_top_in[77], chanx_left_in[19], chanx_left_in[71]}),
		.sram(mux_tree_tapbuf_L1SB_size4_1_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_1_sram_inv[0:1]),
		.out(chanx_right_out[0]));

	mux_tree_tapbuf_L1SB_size4 mux_right_track_36 (
		.in({chany_top_in[17], chany_top_in[56], chany_top_in[95], chanx_left_in[43]}),
		.sram(mux_tree_tapbuf_L1SB_size4_2_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_2_sram_inv[0:1]),
		.out(chanx_right_out[18]));

	mux_tree_tapbuf_L1SB_size4 mux_left_track_3 (
		.in({chany_top_in[38], chany_top_in[77], chanx_right_in[20], chanx_right_in[72]}),
		.sram(mux_tree_tapbuf_L1SB_size4_3_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_3_sram_inv[0:1]),
		.out(chanx_left_out[1]));

	mux_tree_tapbuf_L1SB_size4 mux_left_track_5 (
		.in({chany_top_in[37], chany_top_in[76], chanx_right_in[21], chanx_right_in[73]}),
		.sram(mux_tree_tapbuf_L1SB_size4_4_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_4_sram_inv[0:1]),
		.out(chanx_left_out[2]));

	mux_tree_tapbuf_L1SB_size4 mux_left_track_7 (
		.in({chany_top_in[36], chany_top_in[75], chanx_right_in[23], chanx_right_in[75]}),
		.sram(mux_tree_tapbuf_L1SB_size4_5_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_5_sram_inv[0:1]),
		.out(chanx_left_out[3]));

	mux_tree_tapbuf_L1SB_size4 mux_left_track_9 (
		.in({chany_top_in[35], chany_top_in[74], chanx_right_in[24], chanx_right_in[76]}),
		.sram(mux_tree_tapbuf_L1SB_size4_6_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_6_sram_inv[0:1]),
		.out(chanx_left_out[4]));

	mux_tree_tapbuf_L1SB_size4 mux_left_track_11 (
		.in({chany_top_in[34], chany_top_in[73], chanx_right_in[25], chanx_right_in[77]}),
		.sram(mux_tree_tapbuf_L1SB_size4_7_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_7_sram_inv[0:1]),
		.out(chanx_left_out[5]));

	mux_tree_tapbuf_L1SB_size4 mux_left_track_13 (
		.in({chany_top_in[33], chany_top_in[72], chanx_right_in[27], chanx_right_in[79]}),
		.sram(mux_tree_tapbuf_L1SB_size4_8_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_8_sram_inv[0:1]),
		.out(chanx_left_out[6]));

	mux_tree_tapbuf_L1SB_size4 mux_left_track_15 (
		.in({chany_top_in[32], chany_top_in[71], chanx_right_in[28], chanx_right_in[80]}),
		.sram(mux_tree_tapbuf_L1SB_size4_9_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_9_sram_inv[0:1]),
		.out(chanx_left_out[7]));

	mux_tree_tapbuf_L1SB_size4 mux_left_track_17 (
		.in({chany_top_in[31], chany_top_in[70], chanx_right_in[29], chanx_right_in[81]}),
		.sram(mux_tree_tapbuf_L1SB_size4_10_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_10_sram_inv[0:1]),
		.out(chanx_left_out[8]));

	mux_tree_tapbuf_L1SB_size4 mux_left_track_19 (
		.in({chany_top_in[30], chany_top_in[69], chanx_right_in[31], chanx_right_in[83]}),
		.sram(mux_tree_tapbuf_L1SB_size4_11_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_11_sram_inv[0:1]),
		.out(chanx_left_out[9]));

	mux_tree_tapbuf_L1SB_size4 mux_left_track_21 (
		.in({chany_top_in[29], chany_top_in[68], chanx_right_in[32], chanx_right_in[84]}),
		.sram(mux_tree_tapbuf_L1SB_size4_12_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_12_sram_inv[0:1]),
		.out(chanx_left_out[10]));

	mux_tree_tapbuf_L1SB_size4 mux_left_track_23 (
		.in({chany_top_in[28], chany_top_in[67], chanx_right_in[33], chanx_right_in[85]}),
		.sram(mux_tree_tapbuf_L1SB_size4_13_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_13_sram_inv[0:1]),
		.out(chanx_left_out[11]));

	mux_tree_tapbuf_L1SB_size4 mux_left_track_25 (
		.in({chany_top_in[27], chany_top_in[66], chanx_right_in[35], chanx_right_in[87]}),
		.sram(mux_tree_tapbuf_L1SB_size4_14_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_14_sram_inv[0:1]),
		.out(chanx_left_out[12]));

	mux_tree_tapbuf_L1SB_size4 mux_left_track_27 (
		.in({chany_top_in[26], chany_top_in[65], chanx_right_in[36], chanx_right_in[88]}),
		.sram(mux_tree_tapbuf_L1SB_size4_15_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_15_sram_inv[0:1]),
		.out(chanx_left_out[13]));

	mux_tree_tapbuf_L1SB_size4 mux_left_track_29 (
		.in({chany_top_in[25], chany_top_in[64], chanx_right_in[37], chanx_right_in[89]}),
		.sram(mux_tree_tapbuf_L1SB_size4_16_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_16_sram_inv[0:1]),
		.out(chanx_left_out[14]));

	mux_tree_tapbuf_L1SB_size4 mux_left_track_31 (
		.in({chany_top_in[24], chany_top_in[63], chanx_right_in[39], chanx_right_in[91]}),
		.sram(mux_tree_tapbuf_L1SB_size4_17_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_17_sram_inv[0:1]),
		.out(chanx_left_out[15]));

	mux_tree_tapbuf_L1SB_size4 mux_left_track_33 (
		.in({chany_top_in[23], chany_top_in[62], chanx_right_in[40], chanx_right_in[92]}),
		.sram(mux_tree_tapbuf_L1SB_size4_18_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_18_sram_inv[0:1]),
		.out(chanx_left_out[16]));

	mux_tree_tapbuf_L1SB_size4 mux_left_track_35 (
		.in({chany_top_in[22], chany_top_in[61], chanx_right_in[41], chanx_right_in[93]}),
		.sram(mux_tree_tapbuf_L1SB_size4_19_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size4_19_sram_inv[0:1]),
		.out(chanx_left_out[17]));

	mux_tree_tapbuf_L1SB_size4_mem mem_top_track_0 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(ccff_head),
		.ccff_tail(mux_tree_tapbuf_L1SB_size4_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size4_0_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_0_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size4_mem mem_right_track_0 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size2_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size4_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size4_1_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_1_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size4_mem mem_right_track_36 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size5_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size4_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size4_2_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_2_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size4_mem mem_left_track_3 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size5_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size4_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size4_3_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_3_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size4_mem mem_left_track_5 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size4_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size4_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size4_4_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_4_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size4_mem mem_left_track_7 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size4_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size4_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size4_5_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_5_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size4_mem mem_left_track_9 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size4_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size4_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size4_6_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_6_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size4_mem mem_left_track_11 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size4_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size4_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size4_7_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_7_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size4_mem mem_left_track_13 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size4_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size4_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size4_8_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_8_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size4_mem mem_left_track_15 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size4_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size4_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size4_9_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_9_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size4_mem mem_left_track_17 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size4_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size4_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size4_10_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_10_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size4_mem mem_left_track_19 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size4_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size4_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size4_11_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_11_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size4_mem mem_left_track_21 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size4_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size4_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size4_12_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_12_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size4_mem mem_left_track_23 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size4_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size4_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size4_13_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_13_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size4_mem mem_left_track_25 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size4_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size4_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size4_14_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_14_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size4_mem mem_left_track_27 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size4_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size4_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size4_15_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_15_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size4_mem mem_left_track_29 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size4_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size4_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size4_16_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_16_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size4_mem mem_left_track_31 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size4_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size4_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size4_17_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_17_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size4_mem mem_left_track_33 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size4_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size4_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size4_18_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_18_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size4_mem mem_left_track_35 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size4_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size4_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size4_19_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size4_19_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size3 mux_top_track_2 (
		.in({chanx_right_in[2], chanx_right_in[20], chanx_left_in[20]}),
		.sram(mux_tree_tapbuf_L1SB_size3_0_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size3_0_sram_inv[0:1]),
		.out(chany_top_out[1]));

	mux_tree_tapbuf_L1SB_size3 mux_top_track_4 (
		.in({chanx_right_in[3], chanx_right_in[21], chanx_left_in[21]}),
		.sram(mux_tree_tapbuf_L1SB_size3_1_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size3_1_sram_inv[0:1]),
		.out(chany_top_out[2]));

	mux_tree_tapbuf_L1SB_size3 mux_top_track_6 (
		.in({chanx_right_in[4], chanx_right_in[23], chanx_left_in[23]}),
		.sram(mux_tree_tapbuf_L1SB_size3_2_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size3_2_sram_inv[0:1]),
		.out(chany_top_out[3]));

	mux_tree_tapbuf_L1SB_size3 mux_top_track_8 (
		.in({chanx_right_in[5], chanx_right_in[24], chanx_left_in[24]}),
		.sram(mux_tree_tapbuf_L1SB_size3_3_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size3_3_sram_inv[0:1]),
		.out(chany_top_out[4]));

	mux_tree_tapbuf_L1SB_size3 mux_top_track_10 (
		.in({chanx_right_in[6], chanx_right_in[25], chanx_left_in[25]}),
		.sram(mux_tree_tapbuf_L1SB_size3_4_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size3_4_sram_inv[0:1]),
		.out(chany_top_out[5]));

	mux_tree_tapbuf_L1SB_size3 mux_top_track_12 (
		.in({chanx_right_in[7], chanx_right_in[27], chanx_left_in[27]}),
		.sram(mux_tree_tapbuf_L1SB_size3_5_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size3_5_sram_inv[0:1]),
		.out(chany_top_out[6]));

	mux_tree_tapbuf_L1SB_size3 mux_top_track_14 (
		.in({chanx_right_in[8], chanx_right_in[28], chanx_left_in[28]}),
		.sram(mux_tree_tapbuf_L1SB_size3_6_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size3_6_sram_inv[0:1]),
		.out(chany_top_out[7]));

	mux_tree_tapbuf_L1SB_size3 mux_top_track_16 (
		.in({chanx_right_in[9], chanx_right_in[29], chanx_left_in[29]}),
		.sram(mux_tree_tapbuf_L1SB_size3_7_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size3_7_sram_inv[0:1]),
		.out(chany_top_out[8]));

	mux_tree_tapbuf_L1SB_size3 mux_top_track_18 (
		.in({chanx_right_in[10], chanx_right_in[31], chanx_left_in[31]}),
		.sram(mux_tree_tapbuf_L1SB_size3_8_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size3_8_sram_inv[0:1]),
		.out(chany_top_out[9]));

	mux_tree_tapbuf_L1SB_size3 mux_top_track_20 (
		.in({chanx_right_in[11], chanx_right_in[32], chanx_left_in[32]}),
		.sram(mux_tree_tapbuf_L1SB_size3_9_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size3_9_sram_inv[0:1]),
		.out(chany_top_out[10]));

	mux_tree_tapbuf_L1SB_size3 mux_top_track_22 (
		.in({chanx_right_in[12], chanx_right_in[33], chanx_left_in[33]}),
		.sram(mux_tree_tapbuf_L1SB_size3_10_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size3_10_sram_inv[0:1]),
		.out(chany_top_out[11]));

	mux_tree_tapbuf_L1SB_size3 mux_top_track_24 (
		.in({chanx_right_in[13], chanx_right_in[35], chanx_left_in[35]}),
		.sram(mux_tree_tapbuf_L1SB_size3_11_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size3_11_sram_inv[0:1]),
		.out(chany_top_out[12]));

	mux_tree_tapbuf_L1SB_size3 mux_top_track_26 (
		.in({chanx_right_in[14], chanx_right_in[36], chanx_left_in[36]}),
		.sram(mux_tree_tapbuf_L1SB_size3_12_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size3_12_sram_inv[0:1]),
		.out(chany_top_out[13]));

	mux_tree_tapbuf_L1SB_size3 mux_top_track_28 (
		.in({chanx_right_in[15], chanx_right_in[37], chanx_left_in[37]}),
		.sram(mux_tree_tapbuf_L1SB_size3_13_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size3_13_sram_inv[0:1]),
		.out(chany_top_out[14]));

	mux_tree_tapbuf_L1SB_size3 mux_top_track_30 (
		.in({chanx_right_in[16], chanx_right_in[39], chanx_left_in[39]}),
		.sram(mux_tree_tapbuf_L1SB_size3_14_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size3_14_sram_inv[0:1]),
		.out(chany_top_out[15]));

	mux_tree_tapbuf_L1SB_size3 mux_top_track_32 (
		.in({chanx_right_in[17], chanx_right_in[40], chanx_left_in[40]}),
		.sram(mux_tree_tapbuf_L1SB_size3_15_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size3_15_sram_inv[0:1]),
		.out(chany_top_out[16]));

	mux_tree_tapbuf_L1SB_size3 mux_top_track_34 (
		.in({chanx_right_in[18], chanx_right_in[41], chanx_left_in[41]}),
		.sram(mux_tree_tapbuf_L1SB_size3_16_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size3_16_sram_inv[0:1]),
		.out(chany_top_out[17]));

	mux_tree_tapbuf_L1SB_size3 mux_top_track_36 (
		.in({chanx_right_in[22], chanx_right_in[43], chanx_left_in[43]}),
		.sram(mux_tree_tapbuf_L1SB_size3_17_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size3_17_sram_inv[0:1]),
		.out(chany_top_out[18]));

	mux_tree_tapbuf_L1SB_size3 mux_left_track_37 (
		.in({chany_top_in[21], chany_top_in[60], chanx_right_in[43]}),
		.sram(mux_tree_tapbuf_L1SB_size3_18_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L1SB_size3_18_sram_inv[0:1]),
		.out(chanx_left_out[18]));

	mux_tree_tapbuf_L1SB_size3_mem mem_top_track_2 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size4_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size3_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size3_0_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size3_0_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size3_mem mem_top_track_4 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size3_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size3_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size3_1_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size3_1_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size3_mem mem_top_track_6 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size3_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size3_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size3_2_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size3_2_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size3_mem mem_top_track_8 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size3_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size3_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size3_3_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size3_3_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size3_mem mem_top_track_10 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size3_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size3_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size3_4_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size3_4_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size3_mem mem_top_track_12 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size3_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size3_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size3_5_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size3_5_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size3_mem mem_top_track_14 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size3_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size3_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size3_6_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size3_6_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size3_mem mem_top_track_16 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size3_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size3_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size3_7_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size3_7_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size3_mem mem_top_track_18 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size3_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size3_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size3_8_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size3_8_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size3_mem mem_top_track_20 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size3_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size3_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size3_9_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size3_9_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size3_mem mem_top_track_22 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size3_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size3_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size3_10_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size3_10_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size3_mem mem_top_track_24 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size3_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size3_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size3_11_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size3_11_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size3_mem mem_top_track_26 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size3_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size3_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size3_12_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size3_12_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size3_mem mem_top_track_28 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size3_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size3_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size3_13_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size3_13_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size3_mem mem_top_track_30 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size3_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size3_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size3_14_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size3_14_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size3_mem mem_top_track_32 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size3_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size3_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size3_15_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size3_15_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size3_mem mem_top_track_34 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size3_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size3_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size3_16_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size3_16_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size3_mem mem_top_track_36 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size3_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size3_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size3_17_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size3_17_sram_inv[0:1]));

	mux_tree_tapbuf_L1SB_size3_mem mem_left_track_37 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size4_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size3_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size3_18_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L1SB_size3_18_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3 mux_top_track_38 (
		.in({chanx_right_in[26], chanx_right_in[44], chanx_left_in[44]}),
		.sram(mux_tree_tapbuf_L4SB_size3_0_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_0_sram_inv[0:1]),
		.out(chany_top_out[19]));

	mux_tree_tapbuf_L4SB_size3 mux_top_track_40 (
		.in({chanx_right_in[30], chanx_right_in[45], chanx_left_in[45]}),
		.sram(mux_tree_tapbuf_L4SB_size3_1_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_1_sram_inv[0:1]),
		.out(chany_top_out[20]));

	mux_tree_tapbuf_L4SB_size3 mux_top_track_42 (
		.in({chanx_right_in[34], chanx_right_in[47], chanx_left_in[47]}),
		.sram(mux_tree_tapbuf_L4SB_size3_2_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_2_sram_inv[0:1]),
		.out(chany_top_out[21]));

	mux_tree_tapbuf_L4SB_size3 mux_top_track_44 (
		.in({chanx_right_in[38], chanx_right_in[48], chanx_left_in[48]}),
		.sram(mux_tree_tapbuf_L4SB_size3_3_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_3_sram_inv[0:1]),
		.out(chany_top_out[22]));

	mux_tree_tapbuf_L4SB_size3 mux_top_track_46 (
		.in({chanx_right_in[42], chanx_right_in[49], chanx_left_in[49]}),
		.sram(mux_tree_tapbuf_L4SB_size3_4_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_4_sram_inv[0:1]),
		.out(chany_top_out[23]));

	mux_tree_tapbuf_L4SB_size3 mux_top_track_48 (
		.in({chanx_right_in[46], chanx_right_in[51], chanx_left_in[51]}),
		.sram(mux_tree_tapbuf_L4SB_size3_5_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_5_sram_inv[0:1]),
		.out(chany_top_out[24]));

	mux_tree_tapbuf_L4SB_size3 mux_top_track_50 (
		.in({chanx_right_in[50], chanx_right_in[52], chanx_left_in[52]}),
		.sram(mux_tree_tapbuf_L4SB_size3_6_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_6_sram_inv[0:1]),
		.out(chany_top_out[25]));

	mux_tree_tapbuf_L4SB_size3 mux_top_track_52 (
		.in({chanx_right_in[53:54], chanx_left_in[53]}),
		.sram(mux_tree_tapbuf_L4SB_size3_7_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_7_sram_inv[0:1]),
		.out(chany_top_out[26]));

	mux_tree_tapbuf_L4SB_size3 mux_top_track_54 (
		.in({chanx_right_in[55], chanx_right_in[58], chanx_left_in[55]}),
		.sram(mux_tree_tapbuf_L4SB_size3_8_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_8_sram_inv[0:1]),
		.out(chany_top_out[27]));

	mux_tree_tapbuf_L4SB_size3 mux_top_track_56 (
		.in({chanx_right_in[56], chanx_right_in[62], chanx_left_in[56]}),
		.sram(mux_tree_tapbuf_L4SB_size3_9_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_9_sram_inv[0:1]),
		.out(chany_top_out[28]));

	mux_tree_tapbuf_L4SB_size3 mux_top_track_58 (
		.in({chanx_right_in[57], chanx_right_in[66], chanx_left_in[57]}),
		.sram(mux_tree_tapbuf_L4SB_size3_10_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_10_sram_inv[0:1]),
		.out(chany_top_out[29]));

	mux_tree_tapbuf_L4SB_size3 mux_top_track_60 (
		.in({chanx_right_in[59], chanx_right_in[70], chanx_left_in[59]}),
		.sram(mux_tree_tapbuf_L4SB_size3_11_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_11_sram_inv[0:1]),
		.out(chany_top_out[30]));

	mux_tree_tapbuf_L4SB_size3 mux_top_track_62 (
		.in({chanx_right_in[60], chanx_right_in[74], chanx_left_in[60]}),
		.sram(mux_tree_tapbuf_L4SB_size3_12_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_12_sram_inv[0:1]),
		.out(chany_top_out[31]));

	mux_tree_tapbuf_L4SB_size3 mux_top_track_64 (
		.in({chanx_right_in[61], chanx_right_in[78], chanx_left_in[61]}),
		.sram(mux_tree_tapbuf_L4SB_size3_13_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_13_sram_inv[0:1]),
		.out(chany_top_out[32]));

	mux_tree_tapbuf_L4SB_size3 mux_top_track_66 (
		.in({chanx_right_in[63], chanx_right_in[82], chanx_left_in[63]}),
		.sram(mux_tree_tapbuf_L4SB_size3_14_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_14_sram_inv[0:1]),
		.out(chany_top_out[33]));

	mux_tree_tapbuf_L4SB_size3 mux_top_track_68 (
		.in({chanx_right_in[64], chanx_right_in[86], chanx_left_in[64]}),
		.sram(mux_tree_tapbuf_L4SB_size3_15_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_15_sram_inv[0:1]),
		.out(chany_top_out[34]));

	mux_tree_tapbuf_L4SB_size3 mux_top_track_70 (
		.in({chanx_right_in[65], chanx_right_in[90], chanx_left_in[65]}),
		.sram(mux_tree_tapbuf_L4SB_size3_16_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_16_sram_inv[0:1]),
		.out(chany_top_out[35]));

	mux_tree_tapbuf_L4SB_size3 mux_top_track_72 (
		.in({chanx_right_in[67], chanx_right_in[94], chanx_left_in[67]}),
		.sram(mux_tree_tapbuf_L4SB_size3_17_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_17_sram_inv[0:1]),
		.out(chany_top_out[36]));

	mux_tree_tapbuf_L4SB_size3 mux_top_track_74 (
		.in({chanx_right_in[68], chanx_right_in[95], chanx_left_in[68]}),
		.sram(mux_tree_tapbuf_L4SB_size3_18_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_18_sram_inv[0:1]),
		.out(chany_top_out[37]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_38 (
		.in({chany_top_in[18], chany_top_in[57], chanx_left_in[44]}),
		.sram(mux_tree_tapbuf_L4SB_size3_19_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_19_sram_inv[0:1]),
		.out(chanx_right_out[19]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_46 (
		.in({chany_top_in[19], chany_top_in[58], chanx_left_in[45]}),
		.sram(mux_tree_tapbuf_L4SB_size3_20_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_20_sram_inv[0:1]),
		.out(chanx_right_out[23]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_54 (
		.in({chany_top_in[20], chany_top_in[59], chanx_left_in[47]}),
		.sram(mux_tree_tapbuf_L4SB_size3_21_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_21_sram_inv[0:1]),
		.out(chanx_right_out[27]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_62 (
		.in({chany_top_in[21], chany_top_in[60], chanx_left_in[48]}),
		.sram(mux_tree_tapbuf_L4SB_size3_22_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_22_sram_inv[0:1]),
		.out(chanx_right_out[31]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_70 (
		.in({chany_top_in[22], chany_top_in[61], chanx_left_in[49]}),
		.sram(mux_tree_tapbuf_L4SB_size3_23_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_23_sram_inv[0:1]),
		.out(chanx_right_out[35]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_78 (
		.in({chany_top_in[23], chany_top_in[62], chanx_left_in[51]}),
		.sram(mux_tree_tapbuf_L4SB_size3_24_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_24_sram_inv[0:1]),
		.out(chanx_right_out[39]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_86 (
		.in({chany_top_in[24], chany_top_in[63], chanx_left_in[52]}),
		.sram(mux_tree_tapbuf_L4SB_size3_25_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_25_sram_inv[0:1]),
		.out(chanx_right_out[43]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_94 (
		.in({chany_top_in[25], chany_top_in[64], chanx_left_in[53]}),
		.sram(mux_tree_tapbuf_L4SB_size3_26_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_26_sram_inv[0:1]),
		.out(chanx_right_out[47]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_102 (
		.in({chany_top_in[26], chany_top_in[65], chanx_left_in[55]}),
		.sram(mux_tree_tapbuf_L4SB_size3_27_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_27_sram_inv[0:1]),
		.out(chanx_right_out[51]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_110 (
		.in({chany_top_in[27], chany_top_in[66], chanx_left_in[56]}),
		.sram(mux_tree_tapbuf_L4SB_size3_28_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_28_sram_inv[0:1]),
		.out(chanx_right_out[55]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_118 (
		.in({chany_top_in[28], chany_top_in[67], chanx_left_in[57]}),
		.sram(mux_tree_tapbuf_L4SB_size3_29_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_29_sram_inv[0:1]),
		.out(chanx_right_out[59]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_126 (
		.in({chany_top_in[29], chany_top_in[68], chanx_left_in[59]}),
		.sram(mux_tree_tapbuf_L4SB_size3_30_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_30_sram_inv[0:1]),
		.out(chanx_right_out[63]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_134 (
		.in({chany_top_in[30], chany_top_in[69], chanx_left_in[60]}),
		.sram(mux_tree_tapbuf_L4SB_size3_31_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_31_sram_inv[0:1]),
		.out(chanx_right_out[67]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_142 (
		.in({chany_top_in[31], chany_top_in[70], chanx_left_in[61]}),
		.sram(mux_tree_tapbuf_L4SB_size3_32_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_32_sram_inv[0:1]),
		.out(chanx_right_out[71]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_150 (
		.in({chany_top_in[32], chany_top_in[71], chanx_left_in[63]}),
		.sram(mux_tree_tapbuf_L4SB_size3_33_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_33_sram_inv[0:1]),
		.out(chanx_right_out[75]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_158 (
		.in({chany_top_in[33], chany_top_in[72], chanx_left_in[64]}),
		.sram(mux_tree_tapbuf_L4SB_size3_34_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_34_sram_inv[0:1]),
		.out(chanx_right_out[79]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_166 (
		.in({chany_top_in[34], chany_top_in[73], chanx_left_in[65]}),
		.sram(mux_tree_tapbuf_L4SB_size3_35_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_35_sram_inv[0:1]),
		.out(chanx_right_out[83]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_174 (
		.in({chany_top_in[35], chany_top_in[74], chanx_left_in[67]}),
		.sram(mux_tree_tapbuf_L4SB_size3_36_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_36_sram_inv[0:1]),
		.out(chanx_right_out[87]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_182 (
		.in({chany_top_in[36], chany_top_in[75], chanx_left_in[68]}),
		.sram(mux_tree_tapbuf_L4SB_size3_37_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_37_sram_inv[0:1]),
		.out(chanx_right_out[91]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_190 (
		.in({chany_top_in[37], chany_top_in[76], chanx_left_in[69]}),
		.sram(mux_tree_tapbuf_L4SB_size3_38_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_38_sram_inv[0:1]),
		.out(chanx_right_out[95]));

	mux_tree_tapbuf_L4SB_size3 mux_left_track_39 (
		.in({chany_top_in[20], chany_top_in[59], chanx_right_in[44]}),
		.sram(mux_tree_tapbuf_L4SB_size3_39_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_39_sram_inv[0:1]),
		.out(chanx_left_out[19]));

	mux_tree_tapbuf_L4SB_size3 mux_left_track_47 (
		.in({chany_top_in[19], chany_top_in[58], chanx_right_in[45]}),
		.sram(mux_tree_tapbuf_L4SB_size3_40_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_40_sram_inv[0:1]),
		.out(chanx_left_out[23]));

	mux_tree_tapbuf_L4SB_size3 mux_left_track_55 (
		.in({chany_top_in[18], chany_top_in[57], chanx_right_in[47]}),
		.sram(mux_tree_tapbuf_L4SB_size3_41_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_41_sram_inv[0:1]),
		.out(chanx_left_out[27]));

	mux_tree_tapbuf_L4SB_size3_mem mem_top_track_38 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size3_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_0_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_0_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_top_track_40 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_1_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_1_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_top_track_42 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_2_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_2_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_top_track_44 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_3_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_3_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_top_track_46 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_4_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_4_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_top_track_48 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_5_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_5_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_top_track_50 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_6_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_6_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_top_track_52 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_7_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_7_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_top_track_54 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_8_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_8_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_top_track_56 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_9_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_9_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_top_track_58 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_10_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_10_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_top_track_60 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_11_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_11_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_top_track_62 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_12_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_12_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_top_track_64 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_13_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_13_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_top_track_66 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_14_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_14_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_top_track_68 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_15_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_15_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_top_track_70 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_16_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_16_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_top_track_72 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_17_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_17_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_top_track_74 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_18_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_18_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_38 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size4_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_19_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_19_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_46 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_20_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_20_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_54 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_21_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_21_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_62 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_22_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_22_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_70 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_23_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_23_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_78 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_24_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_24_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_86 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_25_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_25_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_94 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_26_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_26_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_102 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_27_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_27_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_27_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_110 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_27_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_28_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_28_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_28_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_118 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_28_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_29_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_29_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_29_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_126 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_29_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_30_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_30_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_30_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_134 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_30_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_31_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_31_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_31_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_142 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_31_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_32_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_32_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_32_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_150 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_32_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_33_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_33_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_33_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_158 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_33_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_34_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_34_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_34_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_166 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_34_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_35_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_35_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_35_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_174 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_35_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_36_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_36_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_36_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_182 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_36_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_37_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_37_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_37_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_190 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_37_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_38_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_38_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_38_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_left_track_39 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size3_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_39_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_39_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_39_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_left_track_47 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_39_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_40_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_40_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_40_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_left_track_55 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_40_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_41_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_41_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_41_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size2 mux_top_track_76 (
		.in({chanx_right_in[69], chanx_left_in[69]}),
		.sram(mux_tree_tapbuf_L4SB_size2_0_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_0_sram_inv),
		.out(chany_top_out[38]));

	mux_tree_tapbuf_L4SB_size2 mux_top_track_78 (
		.in({chanx_right_in[71], chanx_left_in[71]}),
		.sram(mux_tree_tapbuf_L4SB_size2_1_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_1_sram_inv),
		.out(chany_top_out[39]));

	mux_tree_tapbuf_L4SB_size2 mux_top_track_80 (
		.in({chanx_right_in[72], chanx_left_in[72]}),
		.sram(mux_tree_tapbuf_L4SB_size2_2_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_2_sram_inv),
		.out(chany_top_out[40]));

	mux_tree_tapbuf_L4SB_size2 mux_top_track_82 (
		.in({chanx_right_in[73], chanx_left_in[73]}),
		.sram(mux_tree_tapbuf_L4SB_size2_3_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_3_sram_inv),
		.out(chany_top_out[41]));

	mux_tree_tapbuf_L4SB_size2 mux_top_track_84 (
		.in({chanx_right_in[75], chanx_left_in[75]}),
		.sram(mux_tree_tapbuf_L4SB_size2_4_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_4_sram_inv),
		.out(chany_top_out[42]));

	mux_tree_tapbuf_L4SB_size2 mux_top_track_86 (
		.in({chanx_right_in[76], chanx_left_in[76]}),
		.sram(mux_tree_tapbuf_L4SB_size2_5_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_5_sram_inv),
		.out(chany_top_out[43]));

	mux_tree_tapbuf_L4SB_size2 mux_top_track_88 (
		.in({chanx_right_in[77], chanx_left_in[77]}),
		.sram(mux_tree_tapbuf_L4SB_size2_6_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_6_sram_inv),
		.out(chany_top_out[44]));

	mux_tree_tapbuf_L4SB_size2 mux_top_track_90 (
		.in({chanx_right_in[79], chanx_left_in[79]}),
		.sram(mux_tree_tapbuf_L4SB_size2_7_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_7_sram_inv),
		.out(chany_top_out[45]));

	mux_tree_tapbuf_L4SB_size2 mux_top_track_92 (
		.in({chanx_right_in[80], chanx_left_in[80]}),
		.sram(mux_tree_tapbuf_L4SB_size2_8_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_8_sram_inv),
		.out(chany_top_out[46]));

	mux_tree_tapbuf_L4SB_size2 mux_top_track_94 (
		.in({chanx_right_in[81], chanx_left_in[81]}),
		.sram(mux_tree_tapbuf_L4SB_size2_9_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_9_sram_inv),
		.out(chany_top_out[47]));

	mux_tree_tapbuf_L4SB_size2 mux_top_track_96 (
		.in({chanx_right_in[83], chanx_left_in[83]}),
		.sram(mux_tree_tapbuf_L4SB_size2_10_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_10_sram_inv),
		.out(chany_top_out[48]));

	mux_tree_tapbuf_L4SB_size2 mux_top_track_98 (
		.in({chanx_right_in[84], chanx_left_in[84]}),
		.sram(mux_tree_tapbuf_L4SB_size2_11_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_11_sram_inv),
		.out(chany_top_out[49]));

	mux_tree_tapbuf_L4SB_size2 mux_top_track_100 (
		.in({chanx_right_in[85], chanx_left_in[85]}),
		.sram(mux_tree_tapbuf_L4SB_size2_12_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_12_sram_inv),
		.out(chany_top_out[50]));

	mux_tree_tapbuf_L4SB_size2 mux_top_track_102 (
		.in({chanx_right_in[87], chanx_left_in[87]}),
		.sram(mux_tree_tapbuf_L4SB_size2_13_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_13_sram_inv),
		.out(chany_top_out[51]));

	mux_tree_tapbuf_L4SB_size2 mux_top_track_104 (
		.in({chanx_right_in[88], chanx_left_in[88]}),
		.sram(mux_tree_tapbuf_L4SB_size2_14_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_14_sram_inv),
		.out(chany_top_out[52]));

	mux_tree_tapbuf_L4SB_size2 mux_top_track_106 (
		.in({chanx_right_in[89], chanx_left_in[89]}),
		.sram(mux_tree_tapbuf_L4SB_size2_15_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_15_sram_inv),
		.out(chany_top_out[53]));

	mux_tree_tapbuf_L4SB_size2 mux_top_track_108 (
		.in({chanx_right_in[91], chanx_left_in[91]}),
		.sram(mux_tree_tapbuf_L4SB_size2_16_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_16_sram_inv),
		.out(chany_top_out[54]));

	mux_tree_tapbuf_L4SB_size2 mux_top_track_110 (
		.in({chanx_right_in[92], chanx_left_in[92]}),
		.sram(mux_tree_tapbuf_L4SB_size2_17_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_17_sram_inv),
		.out(chany_top_out[55]));

	mux_tree_tapbuf_L4SB_size2 mux_top_track_112 (
		.in({chanx_right_in[93], chanx_left_in[93]}),
		.sram(mux_tree_tapbuf_L4SB_size2_18_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_18_sram_inv),
		.out(chany_top_out[56]));

	mux_tree_tapbuf_L4SB_size2 mux_top_track_190 (
		.in({chanx_right_in[0], chanx_left_in[1]}),
		.sram(mux_tree_tapbuf_L4SB_size2_19_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_19_sram_inv),
		.out(chany_top_out[95]));

	mux_tree_tapbuf_L4SB_size2_mem mem_top_track_76 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size2_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size2_0_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_0_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_top_track_78 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size2_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size2_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size2_1_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_1_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_top_track_80 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size2_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size2_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size2_2_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_2_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_top_track_82 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size2_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size2_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size2_3_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_3_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_top_track_84 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size2_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size2_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size2_4_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_4_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_top_track_86 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size2_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size2_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size2_5_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_5_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_top_track_88 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size2_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size2_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size2_6_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_6_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_top_track_90 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size2_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size2_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size2_7_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_7_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_top_track_92 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size2_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size2_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size2_8_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_8_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_top_track_94 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size2_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size2_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size2_9_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_9_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_top_track_96 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size2_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size2_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size2_10_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_10_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_top_track_98 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size2_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size2_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size2_11_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_11_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_top_track_100 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size2_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size2_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size2_12_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_12_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_top_track_102 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size2_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size2_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size2_13_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_13_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_top_track_104 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size2_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size2_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size2_14_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_14_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_top_track_106 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size2_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size2_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size2_15_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_15_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_top_track_108 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size2_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size2_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size2_16_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_16_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_top_track_110 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size2_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size2_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size2_17_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_17_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_top_track_112 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size2_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size2_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size2_18_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_18_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_top_track_190 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size2_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size2_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size2_19_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_19_sram_inv));

	mux_tree_tapbuf_L1SB_size5 mux_right_track_2 (
		.in({chany_top_in[0], chany_top_in[39], chany_top_in[78], chanx_left_in[20], chanx_left_in[72]}),
		.sram(mux_tree_tapbuf_L1SB_size5_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size5_0_sram_inv[0:2]),
		.out(chanx_right_out[1]));

	mux_tree_tapbuf_L1SB_size5 mux_right_track_4 (
		.in({chany_top_in[1], chany_top_in[40], chany_top_in[79], chanx_left_in[21], chanx_left_in[73]}),
		.sram(mux_tree_tapbuf_L1SB_size5_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size5_1_sram_inv[0:2]),
		.out(chanx_right_out[2]));

	mux_tree_tapbuf_L1SB_size5 mux_right_track_6 (
		.in({chany_top_in[2], chany_top_in[41], chany_top_in[80], chanx_left_in[23], chanx_left_in[75]}),
		.sram(mux_tree_tapbuf_L1SB_size5_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size5_2_sram_inv[0:2]),
		.out(chanx_right_out[3]));

	mux_tree_tapbuf_L1SB_size5 mux_right_track_8 (
		.in({chany_top_in[3], chany_top_in[42], chany_top_in[81], chanx_left_in[24], chanx_left_in[76]}),
		.sram(mux_tree_tapbuf_L1SB_size5_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size5_3_sram_inv[0:2]),
		.out(chanx_right_out[4]));

	mux_tree_tapbuf_L1SB_size5 mux_right_track_10 (
		.in({chany_top_in[4], chany_top_in[43], chany_top_in[82], chanx_left_in[25], chanx_left_in[77]}),
		.sram(mux_tree_tapbuf_L1SB_size5_4_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size5_4_sram_inv[0:2]),
		.out(chanx_right_out[5]));

	mux_tree_tapbuf_L1SB_size5 mux_right_track_12 (
		.in({chany_top_in[5], chany_top_in[44], chany_top_in[83], chanx_left_in[27], chanx_left_in[79]}),
		.sram(mux_tree_tapbuf_L1SB_size5_5_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size5_5_sram_inv[0:2]),
		.out(chanx_right_out[6]));

	mux_tree_tapbuf_L1SB_size5 mux_right_track_14 (
		.in({chany_top_in[6], chany_top_in[45], chany_top_in[84], chanx_left_in[28], chanx_left_in[80]}),
		.sram(mux_tree_tapbuf_L1SB_size5_6_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size5_6_sram_inv[0:2]),
		.out(chanx_right_out[7]));

	mux_tree_tapbuf_L1SB_size5 mux_right_track_16 (
		.in({chany_top_in[7], chany_top_in[46], chany_top_in[85], chanx_left_in[29], chanx_left_in[81]}),
		.sram(mux_tree_tapbuf_L1SB_size5_7_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size5_7_sram_inv[0:2]),
		.out(chanx_right_out[8]));

	mux_tree_tapbuf_L1SB_size5 mux_right_track_18 (
		.in({chany_top_in[8], chany_top_in[47], chany_top_in[86], chanx_left_in[31], chanx_left_in[83]}),
		.sram(mux_tree_tapbuf_L1SB_size5_8_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size5_8_sram_inv[0:2]),
		.out(chanx_right_out[9]));

	mux_tree_tapbuf_L1SB_size5 mux_right_track_20 (
		.in({chany_top_in[9], chany_top_in[48], chany_top_in[87], chanx_left_in[32], chanx_left_in[84]}),
		.sram(mux_tree_tapbuf_L1SB_size5_9_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size5_9_sram_inv[0:2]),
		.out(chanx_right_out[10]));

	mux_tree_tapbuf_L1SB_size5 mux_right_track_22 (
		.in({chany_top_in[10], chany_top_in[49], chany_top_in[88], chanx_left_in[33], chanx_left_in[85]}),
		.sram(mux_tree_tapbuf_L1SB_size5_10_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size5_10_sram_inv[0:2]),
		.out(chanx_right_out[11]));

	mux_tree_tapbuf_L1SB_size5 mux_right_track_24 (
		.in({chany_top_in[11], chany_top_in[50], chany_top_in[89], chanx_left_in[35], chanx_left_in[87]}),
		.sram(mux_tree_tapbuf_L1SB_size5_11_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size5_11_sram_inv[0:2]),
		.out(chanx_right_out[12]));

	mux_tree_tapbuf_L1SB_size5 mux_right_track_26 (
		.in({chany_top_in[12], chany_top_in[51], chany_top_in[90], chanx_left_in[36], chanx_left_in[88]}),
		.sram(mux_tree_tapbuf_L1SB_size5_12_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size5_12_sram_inv[0:2]),
		.out(chanx_right_out[13]));

	mux_tree_tapbuf_L1SB_size5 mux_right_track_28 (
		.in({chany_top_in[13], chany_top_in[52], chany_top_in[91], chanx_left_in[37], chanx_left_in[89]}),
		.sram(mux_tree_tapbuf_L1SB_size5_13_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size5_13_sram_inv[0:2]),
		.out(chanx_right_out[14]));

	mux_tree_tapbuf_L1SB_size5 mux_right_track_30 (
		.in({chany_top_in[14], chany_top_in[53], chany_top_in[92], chanx_left_in[39], chanx_left_in[91]}),
		.sram(mux_tree_tapbuf_L1SB_size5_14_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size5_14_sram_inv[0:2]),
		.out(chanx_right_out[15]));

	mux_tree_tapbuf_L1SB_size5 mux_right_track_32 (
		.in({chany_top_in[15], chany_top_in[54], chany_top_in[93], chanx_left_in[40], chanx_left_in[92]}),
		.sram(mux_tree_tapbuf_L1SB_size5_15_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size5_15_sram_inv[0:2]),
		.out(chanx_right_out[16]));

	mux_tree_tapbuf_L1SB_size5 mux_right_track_34 (
		.in({chany_top_in[16], chany_top_in[55], chany_top_in[94], chanx_left_in[41], chanx_left_in[93]}),
		.sram(mux_tree_tapbuf_L1SB_size5_16_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size5_16_sram_inv[0:2]),
		.out(chanx_right_out[17]));

	mux_tree_tapbuf_L1SB_size5 mux_left_track_1 (
		.in({chany_top_in[0], chany_top_in[39], chany_top_in[78], chanx_right_in[19], chanx_right_in[71]}),
		.sram(mux_tree_tapbuf_L1SB_size5_17_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size5_17_sram_inv[0:2]),
		.out(chanx_left_out[0]));

	mux_tree_tapbuf_L1SB_size5_mem mem_right_track_2 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size4_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size5_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size5_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size5_0_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size5_mem mem_right_track_4 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size5_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size5_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size5_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size5_1_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size5_mem mem_right_track_6 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size5_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size5_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size5_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size5_2_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size5_mem mem_right_track_8 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size5_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size5_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size5_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size5_3_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size5_mem mem_right_track_10 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size5_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size5_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size5_4_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size5_4_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size5_mem mem_right_track_12 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size5_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size5_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size5_5_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size5_5_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size5_mem mem_right_track_14 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size5_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size5_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size5_6_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size5_6_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size5_mem mem_right_track_16 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size5_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size5_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size5_7_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size5_7_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size5_mem mem_right_track_18 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size5_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size5_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size5_8_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size5_8_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size5_mem mem_right_track_20 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size5_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size5_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size5_9_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size5_9_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size5_mem mem_right_track_22 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size5_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size5_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size5_10_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size5_10_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size5_mem mem_right_track_24 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size5_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size5_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size5_11_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size5_11_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size5_mem mem_right_track_26 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size5_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size5_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size5_12_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size5_12_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size5_mem mem_right_track_28 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size5_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size5_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size5_13_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size5_13_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size5_mem mem_right_track_30 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size5_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size5_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size5_14_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size5_14_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size5_mem mem_right_track_32 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size5_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size5_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size5_15_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size5_15_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size5_mem mem_right_track_34 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size5_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size5_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size5_16_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size5_16_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size5_mem mem_left_track_1 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_38_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size5_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size5_17_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size5_17_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size4 mux_left_track_63 (
		.in({chany_top_in[17], chany_top_in[56], chany_top_in[95], chanx_right_in[48]}),
		.sram(mux_tree_tapbuf_L4SB_size4_0_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_0_sram_inv[0:1]),
		.out(chanx_left_out[31]));

	mux_tree_tapbuf_L4SB_size4 mux_left_track_71 (
		.in({chany_top_in[16], chany_top_in[55], chany_top_in[94], chanx_right_in[49]}),
		.sram(mux_tree_tapbuf_L4SB_size4_1_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_1_sram_inv[0:1]),
		.out(chanx_left_out[35]));

	mux_tree_tapbuf_L4SB_size4 mux_left_track_79 (
		.in({chany_top_in[15], chany_top_in[54], chany_top_in[93], chanx_right_in[51]}),
		.sram(mux_tree_tapbuf_L4SB_size4_2_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_2_sram_inv[0:1]),
		.out(chanx_left_out[39]));

	mux_tree_tapbuf_L4SB_size4 mux_left_track_87 (
		.in({chany_top_in[14], chany_top_in[53], chany_top_in[92], chanx_right_in[52]}),
		.sram(mux_tree_tapbuf_L4SB_size4_3_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_3_sram_inv[0:1]),
		.out(chanx_left_out[43]));

	mux_tree_tapbuf_L4SB_size4 mux_left_track_95 (
		.in({chany_top_in[13], chany_top_in[52], chany_top_in[91], chanx_right_in[53]}),
		.sram(mux_tree_tapbuf_L4SB_size4_4_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_4_sram_inv[0:1]),
		.out(chanx_left_out[47]));

	mux_tree_tapbuf_L4SB_size4 mux_left_track_103 (
		.in({chany_top_in[12], chany_top_in[51], chany_top_in[90], chanx_right_in[55]}),
		.sram(mux_tree_tapbuf_L4SB_size4_5_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_5_sram_inv[0:1]),
		.out(chanx_left_out[51]));

	mux_tree_tapbuf_L4SB_size4 mux_left_track_111 (
		.in({chany_top_in[11], chany_top_in[50], chany_top_in[89], chanx_right_in[56]}),
		.sram(mux_tree_tapbuf_L4SB_size4_6_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_6_sram_inv[0:1]),
		.out(chanx_left_out[55]));

	mux_tree_tapbuf_L4SB_size4 mux_left_track_119 (
		.in({chany_top_in[10], chany_top_in[49], chany_top_in[88], chanx_right_in[57]}),
		.sram(mux_tree_tapbuf_L4SB_size4_7_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_7_sram_inv[0:1]),
		.out(chanx_left_out[59]));

	mux_tree_tapbuf_L4SB_size4 mux_left_track_127 (
		.in({chany_top_in[9], chany_top_in[48], chany_top_in[87], chanx_right_in[59]}),
		.sram(mux_tree_tapbuf_L4SB_size4_8_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_8_sram_inv[0:1]),
		.out(chanx_left_out[63]));

	mux_tree_tapbuf_L4SB_size4 mux_left_track_135 (
		.in({chany_top_in[8], chany_top_in[47], chany_top_in[86], chanx_right_in[60]}),
		.sram(mux_tree_tapbuf_L4SB_size4_9_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_9_sram_inv[0:1]),
		.out(chanx_left_out[67]));

	mux_tree_tapbuf_L4SB_size4 mux_left_track_143 (
		.in({chany_top_in[7], chany_top_in[46], chany_top_in[85], chanx_right_in[61]}),
		.sram(mux_tree_tapbuf_L4SB_size4_10_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_10_sram_inv[0:1]),
		.out(chanx_left_out[71]));

	mux_tree_tapbuf_L4SB_size4 mux_left_track_151 (
		.in({chany_top_in[6], chany_top_in[45], chany_top_in[84], chanx_right_in[63]}),
		.sram(mux_tree_tapbuf_L4SB_size4_11_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_11_sram_inv[0:1]),
		.out(chanx_left_out[75]));

	mux_tree_tapbuf_L4SB_size4 mux_left_track_159 (
		.in({chany_top_in[5], chany_top_in[44], chany_top_in[83], chanx_right_in[64]}),
		.sram(mux_tree_tapbuf_L4SB_size4_12_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_12_sram_inv[0:1]),
		.out(chanx_left_out[79]));

	mux_tree_tapbuf_L4SB_size4 mux_left_track_167 (
		.in({chany_top_in[4], chany_top_in[43], chany_top_in[82], chanx_right_in[65]}),
		.sram(mux_tree_tapbuf_L4SB_size4_13_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_13_sram_inv[0:1]),
		.out(chanx_left_out[83]));

	mux_tree_tapbuf_L4SB_size4 mux_left_track_175 (
		.in({chany_top_in[3], chany_top_in[42], chany_top_in[81], chanx_right_in[67]}),
		.sram(mux_tree_tapbuf_L4SB_size4_14_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_14_sram_inv[0:1]),
		.out(chanx_left_out[87]));

	mux_tree_tapbuf_L4SB_size4 mux_left_track_183 (
		.in({chany_top_in[2], chany_top_in[41], chany_top_in[80], chanx_right_in[68]}),
		.sram(mux_tree_tapbuf_L4SB_size4_15_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_15_sram_inv[0:1]),
		.out(chanx_left_out[91]));

	mux_tree_tapbuf_L4SB_size4 mux_left_track_191 (
		.in({chany_top_in[1], chany_top_in[40], chany_top_in[79], chanx_right_in[69]}),
		.sram(mux_tree_tapbuf_L4SB_size4_16_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size4_16_sram_inv[0:1]),
		.out(chanx_left_out[95]));

	mux_tree_tapbuf_L4SB_size4_mem mem_left_track_63 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_41_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size4_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size4_0_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_0_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_left_track_71 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size4_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size4_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size4_1_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_1_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_left_track_79 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size4_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size4_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size4_2_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_2_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_left_track_87 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size4_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size4_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size4_3_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_3_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_left_track_95 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size4_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size4_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size4_4_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_4_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_left_track_103 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size4_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size4_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size4_5_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_5_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_left_track_111 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size4_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size4_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size4_6_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_6_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_left_track_119 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size4_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size4_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size4_7_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_7_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_left_track_127 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size4_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size4_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size4_8_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_8_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_left_track_135 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size4_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size4_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size4_9_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_9_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_left_track_143 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size4_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size4_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size4_10_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_10_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_left_track_151 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size4_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size4_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size4_11_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_11_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_left_track_159 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size4_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size4_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size4_12_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_12_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_left_track_167 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size4_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size4_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size4_13_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_13_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_left_track_175 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size4_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size4_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size4_14_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_14_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_left_track_183 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size4_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size4_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size4_15_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_15_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size4_mem mem_left_track_191 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size4_mem_15_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size4_16_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size4_16_sram_inv[0:1]));

endmodule
// ----- END Verilog module for sb_2__0_ -----

//----- Default net type -----
`default_nettype none



