//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for Unique Switch Blocks[3][7]
//	Author: Xifan TANG
//	Organization: University of Utah
//-------------------------------------------
//----- Time scale -----
`timescale 1ns / 1ps

//----- Default net type -----
`default_nettype wire

// ----- Verilog module for sb_3__7_ -----
module sb_3__7_(config_enable,
                prog_clock,
                chany_top_in,
                chanx_right_in,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_,
                right_top_grid_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_,
                right_top_grid_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_,
                right_top_grid_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_,
                right_top_grid_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_,
                right_top_grid_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_,
                right_top_grid_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_,
                right_top_grid_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_,
                right_top_grid_bottom_width_0_height_0_subtile_8__pin_a2f_o_0_,
                right_top_grid_bottom_width_0_height_0_subtile_9__pin_a2f_o_0_,
                right_top_grid_bottom_width_0_height_0_subtile_10__pin_a2f_o_0_,
                right_top_grid_bottom_width_0_height_0_subtile_11__pin_a2f_o_0_,
                right_top_grid_bottom_width_0_height_0_subtile_12__pin_a2f_o_0_,
                right_top_grid_bottom_width_0_height_0_subtile_13__pin_a2f_o_0_,
                right_top_grid_bottom_width_0_height_0_subtile_14__pin_a2f_o_0_,
                right_top_grid_bottom_width_0_height_0_subtile_15__pin_a2f_o_0_,
                right_top_grid_bottom_width_0_height_0_subtile_16__pin_a2f_o_0_,
                right_top_grid_bottom_width_0_height_0_subtile_17__pin_a2f_o_0_,
                right_top_grid_bottom_width_0_height_0_subtile_18__pin_a2f_o_0_,
                right_top_grid_bottom_width_0_height_0_subtile_19__pin_a2f_o_0_,
                chany_bottom_in,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_16_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_18_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_19_,
                chanx_left_in,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_,
                left_top_grid_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_,
                left_top_grid_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_,
                left_top_grid_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_,
                left_top_grid_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_,
                left_top_grid_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_,
                left_top_grid_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_,
                left_top_grid_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_,
                left_top_grid_bottom_width_0_height_0_subtile_8__pin_a2f_o_0_,
                left_top_grid_bottom_width_0_height_0_subtile_9__pin_a2f_o_0_,
                left_top_grid_bottom_width_0_height_0_subtile_10__pin_a2f_o_0_,
                left_top_grid_bottom_width_0_height_0_subtile_11__pin_a2f_o_0_,
                left_top_grid_bottom_width_0_height_0_subtile_12__pin_a2f_o_0_,
                left_top_grid_bottom_width_0_height_0_subtile_13__pin_a2f_o_0_,
                left_top_grid_bottom_width_0_height_0_subtile_14__pin_a2f_o_0_,
                left_top_grid_bottom_width_0_height_0_subtile_15__pin_a2f_o_0_,
                left_top_grid_bottom_width_0_height_0_subtile_16__pin_a2f_o_0_,
                left_top_grid_bottom_width_0_height_0_subtile_17__pin_a2f_o_0_,
                left_top_grid_bottom_width_0_height_0_subtile_18__pin_a2f_o_0_,
                left_top_grid_bottom_width_0_height_0_subtile_19__pin_a2f_o_0_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_,
                ccff_head,
                chany_top_out,
                chanx_right_out,
                chany_bottom_out,
                chanx_left_out,
                ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_clock;
//----- INPUT PORTS -----
input [0:95] chany_top_in;
//----- INPUT PORTS -----
input [0:95] chanx_right_in;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_8__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_9__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_10__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_11__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_12__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_13__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_14__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_15__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_16__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_17__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_18__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_19__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:95] chany_bottom_in;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_16_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_18_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_19_;
//----- INPUT PORTS -----
input [0:95] chanx_left_in;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_8__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_9__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_10__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_11__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_12__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_13__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_14__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_15__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_16__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_17__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_18__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_19__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:95] chany_top_out;
//----- OUTPUT PORTS -----
output [0:95] chanx_right_out;
//----- OUTPUT PORTS -----
output [0:95] chany_bottom_out;
//----- OUTPUT PORTS -----
output [0:95] chanx_left_out;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:3] mux_tree_tapbuf_L1SB_size10_0_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size10_0_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size10_10_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size10_10_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size10_11_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size10_11_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size10_1_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size10_1_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size10_2_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size10_2_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size10_3_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size10_3_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size10_4_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size10_4_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size10_5_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size10_5_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size10_6_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size10_6_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size10_7_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size10_7_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size10_8_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size10_8_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size10_9_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size10_9_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size5_0_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size5_0_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size5_1_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size5_1_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size6_0_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size6_0_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size6_1_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size6_1_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size8_0_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size8_0_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size8_10_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size8_10_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size8_11_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size8_11_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size8_12_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size8_12_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size8_13_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size8_13_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size8_14_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size8_14_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size8_15_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size8_15_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size8_16_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size8_16_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size8_17_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size8_17_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size8_18_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size8_18_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size8_19_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size8_19_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size8_1_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size8_1_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size8_20_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size8_20_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size8_21_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size8_21_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size8_22_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size8_22_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size8_23_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size8_23_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size8_24_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size8_24_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size8_25_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size8_25_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size8_2_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size8_2_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size8_3_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size8_3_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size8_4_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size8_4_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size8_5_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size8_5_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size8_6_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size8_6_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size8_7_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size8_7_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size8_8_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size8_8_sram_inv;
wire [0:2] mux_tree_tapbuf_L1SB_size8_9_sram;
wire [0:2] mux_tree_tapbuf_L1SB_size8_9_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_0_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_0_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_10_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_10_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_11_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_11_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_12_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_12_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_13_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_13_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_14_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_14_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_15_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_15_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_16_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_16_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_17_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_17_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_18_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_18_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_19_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_19_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_1_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_1_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_20_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_20_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_21_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_21_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_22_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_22_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_23_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_23_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_24_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_24_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_25_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_25_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_26_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_26_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_27_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_27_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_28_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_28_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_29_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_29_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_2_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_2_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_30_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_30_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_31_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_31_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_32_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_32_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_33_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_33_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_3_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_3_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_4_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_4_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_5_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_5_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_6_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_6_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_7_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_7_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_8_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_8_sram_inv;
wire [0:3] mux_tree_tapbuf_L1SB_size9_9_sram;
wire [0:3] mux_tree_tapbuf_L1SB_size9_9_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size10_0_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size10_0_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size10_1_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size10_1_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size10_2_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size10_2_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size10_3_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size10_3_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size11_0_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size11_0_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size11_10_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size11_10_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size11_11_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size11_11_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size11_1_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size11_1_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size11_2_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size11_2_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size11_3_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size11_3_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size11_4_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size11_4_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size11_5_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size11_5_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size11_6_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size11_6_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size11_7_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size11_7_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size11_8_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size11_8_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size11_9_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size11_9_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size12_0_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size12_0_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size12_1_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size12_1_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size12_2_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size12_2_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size12_3_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size12_3_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_0_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_0_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_10_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_10_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_11_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_11_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_12_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_12_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_13_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_13_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_14_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_14_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_15_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_15_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_16_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_16_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_17_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_17_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_18_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_18_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_19_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_19_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_1_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_1_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_2_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_2_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_3_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_3_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_4_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_4_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_5_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_5_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_6_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_6_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_7_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_7_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_8_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_8_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_9_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_9_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size6_0_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size6_0_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size6_1_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size6_1_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size6_2_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size6_2_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size6_3_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size6_3_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_0_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_0_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_10_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_10_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_11_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_11_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_1_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_1_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_2_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_2_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_3_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_3_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_4_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_4_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_5_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_5_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_6_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_6_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_7_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_7_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_8_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_8_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_9_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_9_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_0_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_0_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_1_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_1_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_2_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_2_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_3_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_3_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_0_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_0_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_10_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_10_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_11_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_11_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_12_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_12_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_13_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_13_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_14_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_14_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_15_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_15_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_16_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_16_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_17_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_17_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_18_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_18_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_19_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_19_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_1_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_1_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_2_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_2_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_3_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_3_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_4_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_4_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_5_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_5_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_6_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_6_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_7_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_7_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_8_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_8_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_9_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_9_sram_inv;

// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 19 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[20] = chany_top_in[19];
// ----- Local connection due to Wire 20 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[21] = chany_top_in[20];
// ----- Local connection due to Wire 21 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[22] = chany_top_in[21];
// ----- Local connection due to Wire 23 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[24] = chany_top_in[23];
// ----- Local connection due to Wire 24 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[25] = chany_top_in[24];
// ----- Local connection due to Wire 25 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[26] = chany_top_in[25];
// ----- Local connection due to Wire 27 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[28] = chany_top_in[27];
// ----- Local connection due to Wire 28 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[29] = chany_top_in[28];
// ----- Local connection due to Wire 29 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[30] = chany_top_in[29];
// ----- Local connection due to Wire 31 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[32] = chany_top_in[31];
// ----- Local connection due to Wire 32 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[33] = chany_top_in[32];
// ----- Local connection due to Wire 33 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[34] = chany_top_in[33];
// ----- Local connection due to Wire 35 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[36] = chany_top_in[35];
// ----- Local connection due to Wire 36 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[37] = chany_top_in[36];
// ----- Local connection due to Wire 37 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[38] = chany_top_in[37];
// ----- Local connection due to Wire 39 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[40] = chany_top_in[39];
// ----- Local connection due to Wire 40 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[41] = chany_top_in[40];
// ----- Local connection due to Wire 41 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[42] = chany_top_in[41];
// ----- Local connection due to Wire 43 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[44] = chany_top_in[43];
// ----- Local connection due to Wire 44 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[45] = chany_top_in[44];
// ----- Local connection due to Wire 45 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[46] = chany_top_in[45];
// ----- Local connection due to Wire 47 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[48] = chany_top_in[47];
// ----- Local connection due to Wire 48 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[49] = chany_top_in[48];
// ----- Local connection due to Wire 49 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[50] = chany_top_in[49];
// ----- Local connection due to Wire 51 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[52] = chany_top_in[51];
// ----- Local connection due to Wire 52 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[53] = chany_top_in[52];
// ----- Local connection due to Wire 53 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[54] = chany_top_in[53];
// ----- Local connection due to Wire 55 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[56] = chany_top_in[55];
// ----- Local connection due to Wire 56 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[57] = chany_top_in[56];
// ----- Local connection due to Wire 57 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[58] = chany_top_in[57];
// ----- Local connection due to Wire 59 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[60] = chany_top_in[59];
// ----- Local connection due to Wire 60 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[61] = chany_top_in[60];
// ----- Local connection due to Wire 61 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[62] = chany_top_in[61];
// ----- Local connection due to Wire 63 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[64] = chany_top_in[63];
// ----- Local connection due to Wire 64 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[65] = chany_top_in[64];
// ----- Local connection due to Wire 65 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[66] = chany_top_in[65];
// ----- Local connection due to Wire 67 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[68] = chany_top_in[67];
// ----- Local connection due to Wire 68 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[69] = chany_top_in[68];
// ----- Local connection due to Wire 69 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[70] = chany_top_in[69];
// ----- Local connection due to Wire 71 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[72] = chany_top_in[71];
// ----- Local connection due to Wire 72 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[73] = chany_top_in[72];
// ----- Local connection due to Wire 73 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[74] = chany_top_in[73];
// ----- Local connection due to Wire 75 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[76] = chany_top_in[75];
// ----- Local connection due to Wire 76 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[77] = chany_top_in[76];
// ----- Local connection due to Wire 77 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[78] = chany_top_in[77];
// ----- Local connection due to Wire 79 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[80] = chany_top_in[79];
// ----- Local connection due to Wire 80 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[81] = chany_top_in[80];
// ----- Local connection due to Wire 81 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[82] = chany_top_in[81];
// ----- Local connection due to Wire 83 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[84] = chany_top_in[83];
// ----- Local connection due to Wire 84 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[85] = chany_top_in[84];
// ----- Local connection due to Wire 85 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[86] = chany_top_in[85];
// ----- Local connection due to Wire 87 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[88] = chany_top_in[87];
// ----- Local connection due to Wire 88 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[89] = chany_top_in[88];
// ----- Local connection due to Wire 89 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[90] = chany_top_in[89];
// ----- Local connection due to Wire 91 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[92] = chany_top_in[91];
// ----- Local connection due to Wire 92 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[93] = chany_top_in[92];
// ----- Local connection due to Wire 93 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_bottom_out[94] = chany_top_in[93];
// ----- Local connection due to Wire 115 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[20] = chanx_right_in[19];
// ----- Local connection due to Wire 116 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[21] = chanx_right_in[20];
// ----- Local connection due to Wire 117 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[22] = chanx_right_in[21];
// ----- Local connection due to Wire 119 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[24] = chanx_right_in[23];
// ----- Local connection due to Wire 120 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[25] = chanx_right_in[24];
// ----- Local connection due to Wire 121 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[26] = chanx_right_in[25];
// ----- Local connection due to Wire 123 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[28] = chanx_right_in[27];
// ----- Local connection due to Wire 124 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[29] = chanx_right_in[28];
// ----- Local connection due to Wire 125 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[30] = chanx_right_in[29];
// ----- Local connection due to Wire 127 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[32] = chanx_right_in[31];
// ----- Local connection due to Wire 128 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[33] = chanx_right_in[32];
// ----- Local connection due to Wire 129 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[34] = chanx_right_in[33];
// ----- Local connection due to Wire 131 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[36] = chanx_right_in[35];
// ----- Local connection due to Wire 132 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[37] = chanx_right_in[36];
// ----- Local connection due to Wire 133 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[38] = chanx_right_in[37];
// ----- Local connection due to Wire 135 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[40] = chanx_right_in[39];
// ----- Local connection due to Wire 136 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[41] = chanx_right_in[40];
// ----- Local connection due to Wire 137 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[42] = chanx_right_in[41];
// ----- Local connection due to Wire 139 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[44] = chanx_right_in[43];
// ----- Local connection due to Wire 140 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[45] = chanx_right_in[44];
// ----- Local connection due to Wire 141 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[46] = chanx_right_in[45];
// ----- Local connection due to Wire 143 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[48] = chanx_right_in[47];
// ----- Local connection due to Wire 144 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[49] = chanx_right_in[48];
// ----- Local connection due to Wire 145 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[50] = chanx_right_in[49];
// ----- Local connection due to Wire 147 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[52] = chanx_right_in[51];
// ----- Local connection due to Wire 148 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[53] = chanx_right_in[52];
// ----- Local connection due to Wire 149 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[54] = chanx_right_in[53];
// ----- Local connection due to Wire 151 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[56] = chanx_right_in[55];
// ----- Local connection due to Wire 152 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[57] = chanx_right_in[56];
// ----- Local connection due to Wire 153 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[58] = chanx_right_in[57];
// ----- Local connection due to Wire 155 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[60] = chanx_right_in[59];
// ----- Local connection due to Wire 156 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[61] = chanx_right_in[60];
// ----- Local connection due to Wire 157 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[62] = chanx_right_in[61];
// ----- Local connection due to Wire 159 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[64] = chanx_right_in[63];
// ----- Local connection due to Wire 160 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[65] = chanx_right_in[64];
// ----- Local connection due to Wire 161 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[66] = chanx_right_in[65];
// ----- Local connection due to Wire 163 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[68] = chanx_right_in[67];
// ----- Local connection due to Wire 164 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[69] = chanx_right_in[68];
// ----- Local connection due to Wire 165 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[70] = chanx_right_in[69];
// ----- Local connection due to Wire 167 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[72] = chanx_right_in[71];
// ----- Local connection due to Wire 168 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[73] = chanx_right_in[72];
// ----- Local connection due to Wire 169 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[74] = chanx_right_in[73];
// ----- Local connection due to Wire 171 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[76] = chanx_right_in[75];
// ----- Local connection due to Wire 172 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[77] = chanx_right_in[76];
// ----- Local connection due to Wire 173 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[78] = chanx_right_in[77];
// ----- Local connection due to Wire 175 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[80] = chanx_right_in[79];
// ----- Local connection due to Wire 176 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[81] = chanx_right_in[80];
// ----- Local connection due to Wire 177 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[82] = chanx_right_in[81];
// ----- Local connection due to Wire 179 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[84] = chanx_right_in[83];
// ----- Local connection due to Wire 180 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[85] = chanx_right_in[84];
// ----- Local connection due to Wire 181 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[86] = chanx_right_in[85];
// ----- Local connection due to Wire 183 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[88] = chanx_right_in[87];
// ----- Local connection due to Wire 184 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[89] = chanx_right_in[88];
// ----- Local connection due to Wire 185 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[90] = chanx_right_in[89];
// ----- Local connection due to Wire 187 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[92] = chanx_right_in[91];
// ----- Local connection due to Wire 188 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[93] = chanx_right_in[92];
// ----- Local connection due to Wire 189 -----
// ----- Net source id 0 -----
// ----- Net sink id 3 -----
	assign chanx_left_out[94] = chanx_right_in[93];
// ----- Local connection due to Wire 231 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[20] = chany_bottom_in[19];
// ----- Local connection due to Wire 232 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[21] = chany_bottom_in[20];
// ----- Local connection due to Wire 233 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[22] = chany_bottom_in[21];
// ----- Local connection due to Wire 235 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[24] = chany_bottom_in[23];
// ----- Local connection due to Wire 236 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[25] = chany_bottom_in[24];
// ----- Local connection due to Wire 237 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[26] = chany_bottom_in[25];
// ----- Local connection due to Wire 239 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[28] = chany_bottom_in[27];
// ----- Local connection due to Wire 240 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[29] = chany_bottom_in[28];
// ----- Local connection due to Wire 241 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[30] = chany_bottom_in[29];
// ----- Local connection due to Wire 243 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[32] = chany_bottom_in[31];
// ----- Local connection due to Wire 244 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[33] = chany_bottom_in[32];
// ----- Local connection due to Wire 245 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[34] = chany_bottom_in[33];
// ----- Local connection due to Wire 247 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[36] = chany_bottom_in[35];
// ----- Local connection due to Wire 248 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[37] = chany_bottom_in[36];
// ----- Local connection due to Wire 249 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[38] = chany_bottom_in[37];
// ----- Local connection due to Wire 251 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[40] = chany_bottom_in[39];
// ----- Local connection due to Wire 252 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[41] = chany_bottom_in[40];
// ----- Local connection due to Wire 253 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[42] = chany_bottom_in[41];
// ----- Local connection due to Wire 255 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[44] = chany_bottom_in[43];
// ----- Local connection due to Wire 256 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[45] = chany_bottom_in[44];
// ----- Local connection due to Wire 257 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[46] = chany_bottom_in[45];
// ----- Local connection due to Wire 259 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[48] = chany_bottom_in[47];
// ----- Local connection due to Wire 260 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[49] = chany_bottom_in[48];
// ----- Local connection due to Wire 261 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[50] = chany_bottom_in[49];
// ----- Local connection due to Wire 263 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[52] = chany_bottom_in[51];
// ----- Local connection due to Wire 264 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[53] = chany_bottom_in[52];
// ----- Local connection due to Wire 265 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[54] = chany_bottom_in[53];
// ----- Local connection due to Wire 267 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[56] = chany_bottom_in[55];
// ----- Local connection due to Wire 268 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[57] = chany_bottom_in[56];
// ----- Local connection due to Wire 269 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[58] = chany_bottom_in[57];
// ----- Local connection due to Wire 271 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[60] = chany_bottom_in[59];
// ----- Local connection due to Wire 272 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[61] = chany_bottom_in[60];
// ----- Local connection due to Wire 273 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[62] = chany_bottom_in[61];
// ----- Local connection due to Wire 275 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[64] = chany_bottom_in[63];
// ----- Local connection due to Wire 276 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[65] = chany_bottom_in[64];
// ----- Local connection due to Wire 277 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[66] = chany_bottom_in[65];
// ----- Local connection due to Wire 279 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[68] = chany_bottom_in[67];
// ----- Local connection due to Wire 280 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[69] = chany_bottom_in[68];
// ----- Local connection due to Wire 281 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[70] = chany_bottom_in[69];
// ----- Local connection due to Wire 283 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[72] = chany_bottom_in[71];
// ----- Local connection due to Wire 284 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[73] = chany_bottom_in[72];
// ----- Local connection due to Wire 285 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[74] = chany_bottom_in[73];
// ----- Local connection due to Wire 287 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[76] = chany_bottom_in[75];
// ----- Local connection due to Wire 288 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[77] = chany_bottom_in[76];
// ----- Local connection due to Wire 289 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[78] = chany_bottom_in[77];
// ----- Local connection due to Wire 291 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[80] = chany_bottom_in[79];
// ----- Local connection due to Wire 292 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[81] = chany_bottom_in[80];
// ----- Local connection due to Wire 293 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[82] = chany_bottom_in[81];
// ----- Local connection due to Wire 295 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[84] = chany_bottom_in[83];
// ----- Local connection due to Wire 296 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[85] = chany_bottom_in[84];
// ----- Local connection due to Wire 297 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[86] = chany_bottom_in[85];
// ----- Local connection due to Wire 299 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[88] = chany_bottom_in[87];
// ----- Local connection due to Wire 300 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[89] = chany_bottom_in[88];
// ----- Local connection due to Wire 301 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[90] = chany_bottom_in[89];
// ----- Local connection due to Wire 303 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[92] = chany_bottom_in[91];
// ----- Local connection due to Wire 304 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[93] = chany_bottom_in[92];
// ----- Local connection due to Wire 305 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_top_out[94] = chany_bottom_in[93];
// ----- Local connection due to Wire 337 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[20] = chanx_left_in[19];
// ----- Local connection due to Wire 338 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[21] = chanx_left_in[20];
// ----- Local connection due to Wire 339 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[22] = chanx_left_in[21];
// ----- Local connection due to Wire 341 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[24] = chanx_left_in[23];
// ----- Local connection due to Wire 342 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[25] = chanx_left_in[24];
// ----- Local connection due to Wire 343 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[26] = chanx_left_in[25];
// ----- Local connection due to Wire 345 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[28] = chanx_left_in[27];
// ----- Local connection due to Wire 346 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[29] = chanx_left_in[28];
// ----- Local connection due to Wire 347 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[30] = chanx_left_in[29];
// ----- Local connection due to Wire 349 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[32] = chanx_left_in[31];
// ----- Local connection due to Wire 350 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[33] = chanx_left_in[32];
// ----- Local connection due to Wire 351 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[34] = chanx_left_in[33];
// ----- Local connection due to Wire 353 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[36] = chanx_left_in[35];
// ----- Local connection due to Wire 354 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[37] = chanx_left_in[36];
// ----- Local connection due to Wire 355 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[38] = chanx_left_in[37];
// ----- Local connection due to Wire 357 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[40] = chanx_left_in[39];
// ----- Local connection due to Wire 358 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[41] = chanx_left_in[40];
// ----- Local connection due to Wire 359 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[42] = chanx_left_in[41];
// ----- Local connection due to Wire 361 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[44] = chanx_left_in[43];
// ----- Local connection due to Wire 362 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[45] = chanx_left_in[44];
// ----- Local connection due to Wire 363 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[46] = chanx_left_in[45];
// ----- Local connection due to Wire 365 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[48] = chanx_left_in[47];
// ----- Local connection due to Wire 366 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[49] = chanx_left_in[48];
// ----- Local connection due to Wire 367 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[50] = chanx_left_in[49];
// ----- Local connection due to Wire 369 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[52] = chanx_left_in[51];
// ----- Local connection due to Wire 370 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[53] = chanx_left_in[52];
// ----- Local connection due to Wire 371 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[54] = chanx_left_in[53];
// ----- Local connection due to Wire 373 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[56] = chanx_left_in[55];
// ----- Local connection due to Wire 374 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[57] = chanx_left_in[56];
// ----- Local connection due to Wire 375 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[58] = chanx_left_in[57];
// ----- Local connection due to Wire 377 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[60] = chanx_left_in[59];
// ----- Local connection due to Wire 378 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[61] = chanx_left_in[60];
// ----- Local connection due to Wire 379 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[62] = chanx_left_in[61];
// ----- Local connection due to Wire 381 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[64] = chanx_left_in[63];
// ----- Local connection due to Wire 382 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[65] = chanx_left_in[64];
// ----- Local connection due to Wire 383 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[66] = chanx_left_in[65];
// ----- Local connection due to Wire 385 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[68] = chanx_left_in[67];
// ----- Local connection due to Wire 386 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[69] = chanx_left_in[68];
// ----- Local connection due to Wire 387 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[70] = chanx_left_in[69];
// ----- Local connection due to Wire 389 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[72] = chanx_left_in[71];
// ----- Local connection due to Wire 390 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[73] = chanx_left_in[72];
// ----- Local connection due to Wire 391 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[74] = chanx_left_in[73];
// ----- Local connection due to Wire 393 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[76] = chanx_left_in[75];
// ----- Local connection due to Wire 394 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[77] = chanx_left_in[76];
// ----- Local connection due to Wire 395 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[78] = chanx_left_in[77];
// ----- Local connection due to Wire 397 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[80] = chanx_left_in[79];
// ----- Local connection due to Wire 398 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[81] = chanx_left_in[80];
// ----- Local connection due to Wire 399 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[82] = chanx_left_in[81];
// ----- Local connection due to Wire 401 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[84] = chanx_left_in[83];
// ----- Local connection due to Wire 402 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[85] = chanx_left_in[84];
// ----- Local connection due to Wire 403 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[86] = chanx_left_in[85];
// ----- Local connection due to Wire 405 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[88] = chanx_left_in[87];
// ----- Local connection due to Wire 406 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[89] = chanx_left_in[88];
// ----- Local connection due to Wire 407 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[90] = chanx_left_in[89];
// ----- Local connection due to Wire 409 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[92] = chanx_left_in[91];
// ----- Local connection due to Wire 410 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[93] = chanx_left_in[92];
// ----- Local connection due to Wire 411 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_right_out[94] = chanx_left_in[93];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	mux_tree_tapbuf_L1SB_size8 mux_top_track_0 (
		.in({chanx_right_in[1], chanx_right_in[19], chanx_right_in[71], chany_bottom_in[19], chany_bottom_in[71], chanx_left_in[0], chanx_left_in[19], chanx_left_in[71]}),
		.sram(mux_tree_tapbuf_L1SB_size8_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size8_0_sram_inv[0:2]),
		.out(chany_top_out[0]));

	mux_tree_tapbuf_L1SB_size8 mux_top_track_2 (
		.in({chanx_right_in[2], chanx_right_in[20], chanx_right_in[72], chany_bottom_in[20], chany_bottom_in[72], chanx_left_in[20], chanx_left_in[72], chanx_left_in[95]}),
		.sram(mux_tree_tapbuf_L1SB_size8_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size8_1_sram_inv[0:2]),
		.out(chany_top_out[1]));

	mux_tree_tapbuf_L1SB_size8 mux_top_track_4 (
		.in({chanx_right_in[3], chanx_right_in[21], chanx_right_in[73], chany_bottom_in[21], chany_bottom_in[73], chanx_left_in[21], chanx_left_in[73], chanx_left_in[94]}),
		.sram(mux_tree_tapbuf_L1SB_size8_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size8_2_sram_inv[0:2]),
		.out(chany_top_out[2]));

	mux_tree_tapbuf_L1SB_size8 mux_top_track_6 (
		.in({chanx_right_in[4], chanx_right_in[23], chanx_right_in[75], chany_bottom_in[23], chany_bottom_in[75], chanx_left_in[23], chanx_left_in[75], chanx_left_in[90]}),
		.sram(mux_tree_tapbuf_L1SB_size8_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size8_3_sram_inv[0:2]),
		.out(chany_top_out[3]));

	mux_tree_tapbuf_L1SB_size8 mux_top_track_8 (
		.in({chanx_right_in[5], chanx_right_in[24], chanx_right_in[76], chany_bottom_in[24], chany_bottom_in[76], chanx_left_in[24], chanx_left_in[76], chanx_left_in[86]}),
		.sram(mux_tree_tapbuf_L1SB_size8_4_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size8_4_sram_inv[0:2]),
		.out(chany_top_out[4]));

	mux_tree_tapbuf_L1SB_size8 mux_top_track_10 (
		.in({chanx_right_in[6], chanx_right_in[25], chanx_right_in[77], chany_bottom_in[25], chany_bottom_in[77], chanx_left_in[25], chanx_left_in[77], chanx_left_in[82]}),
		.sram(mux_tree_tapbuf_L1SB_size8_5_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size8_5_sram_inv[0:2]),
		.out(chany_top_out[5]));

	mux_tree_tapbuf_L1SB_size8 mux_top_track_12 (
		.in({chanx_right_in[7], chanx_right_in[27], chanx_right_in[79], chany_bottom_in[27], chany_bottom_in[79], chanx_left_in[27], chanx_left_in[78:79]}),
		.sram(mux_tree_tapbuf_L1SB_size8_6_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size8_6_sram_inv[0:2]),
		.out(chany_top_out[6]));

	mux_tree_tapbuf_L1SB_size8 mux_top_track_14 (
		.in({chanx_right_in[8], chanx_right_in[28], chanx_right_in[80], chany_bottom_in[28], chany_bottom_in[80], chanx_left_in[28], chanx_left_in[74], chanx_left_in[80]}),
		.sram(mux_tree_tapbuf_L1SB_size8_7_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size8_7_sram_inv[0:2]),
		.out(chany_top_out[7]));

	mux_tree_tapbuf_L1SB_size8 mux_top_track_16 (
		.in({chanx_right_in[9], chanx_right_in[29], chanx_right_in[81], chany_bottom_in[29], chany_bottom_in[81], chanx_left_in[29], chanx_left_in[70], chanx_left_in[81]}),
		.sram(mux_tree_tapbuf_L1SB_size8_8_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size8_8_sram_inv[0:2]),
		.out(chany_top_out[8]));

	mux_tree_tapbuf_L1SB_size8 mux_top_track_18 (
		.in({chanx_right_in[10], chanx_right_in[31], chanx_right_in[83], chany_bottom_in[31], chany_bottom_in[83], chanx_left_in[31], chanx_left_in[66], chanx_left_in[83]}),
		.sram(mux_tree_tapbuf_L1SB_size8_9_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size8_9_sram_inv[0:2]),
		.out(chany_top_out[9]));

	mux_tree_tapbuf_L1SB_size8 mux_top_track_20 (
		.in({chanx_right_in[11], chanx_right_in[32], chanx_right_in[84], chany_bottom_in[32], chany_bottom_in[84], chanx_left_in[32], chanx_left_in[62], chanx_left_in[84]}),
		.sram(mux_tree_tapbuf_L1SB_size8_10_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size8_10_sram_inv[0:2]),
		.out(chany_top_out[10]));

	mux_tree_tapbuf_L1SB_size8 mux_top_track_22 (
		.in({chanx_right_in[12], chanx_right_in[33], chanx_right_in[85], chany_bottom_in[33], chany_bottom_in[85], chanx_left_in[33], chanx_left_in[58], chanx_left_in[85]}),
		.sram(mux_tree_tapbuf_L1SB_size8_11_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size8_11_sram_inv[0:2]),
		.out(chany_top_out[11]));

	mux_tree_tapbuf_L1SB_size8 mux_top_track_24 (
		.in({chanx_right_in[13], chanx_right_in[35], chanx_right_in[87], chany_bottom_in[35], chany_bottom_in[87], chanx_left_in[35], chanx_left_in[54], chanx_left_in[87]}),
		.sram(mux_tree_tapbuf_L1SB_size8_12_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size8_12_sram_inv[0:2]),
		.out(chany_top_out[12]));

	mux_tree_tapbuf_L1SB_size8 mux_top_track_26 (
		.in({chanx_right_in[14], chanx_right_in[36], chanx_right_in[88], chany_bottom_in[36], chany_bottom_in[88], chanx_left_in[36], chanx_left_in[50], chanx_left_in[88]}),
		.sram(mux_tree_tapbuf_L1SB_size8_13_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size8_13_sram_inv[0:2]),
		.out(chany_top_out[13]));

	mux_tree_tapbuf_L1SB_size8 mux_top_track_28 (
		.in({chanx_right_in[15], chanx_right_in[37], chanx_right_in[89], chany_bottom_in[37], chany_bottom_in[89], chanx_left_in[37], chanx_left_in[46], chanx_left_in[89]}),
		.sram(mux_tree_tapbuf_L1SB_size8_14_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size8_14_sram_inv[0:2]),
		.out(chany_top_out[14]));

	mux_tree_tapbuf_L1SB_size8 mux_top_track_30 (
		.in({chanx_right_in[16], chanx_right_in[39], chanx_right_in[91], chany_bottom_in[39], chany_bottom_in[91], chanx_left_in[39], chanx_left_in[42], chanx_left_in[91]}),
		.sram(mux_tree_tapbuf_L1SB_size8_15_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size8_15_sram_inv[0:2]),
		.out(chany_top_out[15]));

	mux_tree_tapbuf_L1SB_size8 mux_top_track_32 (
		.in({chanx_right_in[17], chanx_right_in[40], chanx_right_in[92], chany_bottom_in[40], chany_bottom_in[92], chanx_left_in[38], chanx_left_in[40], chanx_left_in[92]}),
		.sram(mux_tree_tapbuf_L1SB_size8_16_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size8_16_sram_inv[0:2]),
		.out(chany_top_out[16]));

	mux_tree_tapbuf_L1SB_size8 mux_top_track_34 (
		.in({chanx_right_in[18], chanx_right_in[41], chanx_right_in[93], chany_bottom_in[41], chany_bottom_in[93], chanx_left_in[34], chanx_left_in[41], chanx_left_in[93]}),
		.sram(mux_tree_tapbuf_L1SB_size8_17_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size8_17_sram_inv[0:2]),
		.out(chany_top_out[17]));

	mux_tree_tapbuf_L1SB_size8 mux_bottom_track_21 (
		.in({chany_top_in[32], chany_top_in[84], chanx_right_in[32], chanx_right_in[54], chanx_right_in[84], chanx_left_in[11], chanx_left_in[32], chanx_left_in[84]}),
		.sram(mux_tree_tapbuf_L1SB_size8_18_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size8_18_sram_inv[0:2]),
		.out(chany_bottom_out[10]));

	mux_tree_tapbuf_L1SB_size8 mux_bottom_track_23 (
		.in({chany_top_in[33], chany_top_in[85], chanx_right_in[33], chanx_right_in[50], chanx_right_in[85], chanx_left_in[12], chanx_left_in[33], chanx_left_in[85]}),
		.sram(mux_tree_tapbuf_L1SB_size8_19_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size8_19_sram_inv[0:2]),
		.out(chany_bottom_out[11]));

	mux_tree_tapbuf_L1SB_size8 mux_bottom_track_25 (
		.in({chany_top_in[35], chany_top_in[87], chanx_right_in[35], chanx_right_in[46], chanx_right_in[87], chanx_left_in[13], chanx_left_in[35], chanx_left_in[87]}),
		.sram(mux_tree_tapbuf_L1SB_size8_20_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size8_20_sram_inv[0:2]),
		.out(chany_bottom_out[12]));

	mux_tree_tapbuf_L1SB_size8 mux_bottom_track_27 (
		.in({chany_top_in[36], chany_top_in[88], chanx_right_in[36], chanx_right_in[42], chanx_right_in[88], chanx_left_in[14], chanx_left_in[36], chanx_left_in[88]}),
		.sram(mux_tree_tapbuf_L1SB_size8_21_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size8_21_sram_inv[0:2]),
		.out(chany_bottom_out[13]));

	mux_tree_tapbuf_L1SB_size8 mux_bottom_track_29 (
		.in({chany_top_in[37], chany_top_in[89], chanx_right_in[37:38], chanx_right_in[89], chanx_left_in[15], chanx_left_in[37], chanx_left_in[89]}),
		.sram(mux_tree_tapbuf_L1SB_size8_22_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size8_22_sram_inv[0:2]),
		.out(chany_bottom_out[14]));

	mux_tree_tapbuf_L1SB_size8 mux_bottom_track_31 (
		.in({chany_top_in[39], chany_top_in[91], chanx_right_in[34], chanx_right_in[39], chanx_right_in[91], chanx_left_in[16], chanx_left_in[39], chanx_left_in[91]}),
		.sram(mux_tree_tapbuf_L1SB_size8_23_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size8_23_sram_inv[0:2]),
		.out(chany_bottom_out[15]));

	mux_tree_tapbuf_L1SB_size8 mux_bottom_track_33 (
		.in({chany_top_in[40], chany_top_in[92], chanx_right_in[30], chanx_right_in[40], chanx_right_in[92], chanx_left_in[17], chanx_left_in[40], chanx_left_in[92]}),
		.sram(mux_tree_tapbuf_L1SB_size8_24_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size8_24_sram_inv[0:2]),
		.out(chany_bottom_out[16]));

	mux_tree_tapbuf_L1SB_size8 mux_bottom_track_35 (
		.in({chany_top_in[41], chany_top_in[93], chanx_right_in[26], chanx_right_in[41], chanx_right_in[93], chanx_left_in[18], chanx_left_in[41], chanx_left_in[93]}),
		.sram(mux_tree_tapbuf_L1SB_size8_25_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size8_25_sram_inv[0:2]),
		.out(chany_bottom_out[17]));

	mux_tree_tapbuf_L1SB_size8_mem mem_top_track_0 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(ccff_head),
		.ccff_tail(mux_tree_tapbuf_L1SB_size8_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size8_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size8_0_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size8_mem mem_top_track_2 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size8_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size8_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size8_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size8_1_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size8_mem mem_top_track_4 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size8_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size8_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size8_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size8_2_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size8_mem mem_top_track_6 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size8_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size8_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size8_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size8_3_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size8_mem mem_top_track_8 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size8_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size8_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size8_4_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size8_4_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size8_mem mem_top_track_10 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size8_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size8_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size8_5_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size8_5_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size8_mem mem_top_track_12 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size8_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size8_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size8_6_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size8_6_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size8_mem mem_top_track_14 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size8_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size8_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size8_7_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size8_7_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size8_mem mem_top_track_16 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size8_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size8_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size8_8_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size8_8_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size8_mem mem_top_track_18 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size8_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size8_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size8_9_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size8_9_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size8_mem mem_top_track_20 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size8_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size8_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size8_10_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size8_10_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size8_mem mem_top_track_22 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size8_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size8_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size8_11_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size8_11_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size8_mem mem_top_track_24 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size8_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size8_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size8_12_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size8_12_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size8_mem mem_top_track_26 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size8_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size8_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size8_13_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size8_13_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size8_mem mem_top_track_28 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size8_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size8_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size8_14_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size8_14_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size8_mem mem_top_track_30 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size8_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size8_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size8_15_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size8_15_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size8_mem mem_top_track_32 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size8_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size8_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size8_16_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size8_16_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size8_mem mem_top_track_34 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size8_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size8_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size8_17_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size8_17_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size8_mem mem_bottom_track_21 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size9_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size8_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size8_18_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size8_18_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size8_mem mem_bottom_track_23 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size8_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size8_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size8_19_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size8_19_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size8_mem mem_bottom_track_25 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size8_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size8_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size8_20_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size8_20_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size8_mem mem_bottom_track_27 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size8_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size8_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size8_21_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size8_21_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size8_mem mem_bottom_track_29 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size8_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size8_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size8_22_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size8_22_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size8_mem mem_bottom_track_31 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size8_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size8_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size8_23_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size8_23_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size8_mem mem_bottom_track_33 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size8_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size8_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size8_24_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size8_24_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size8_mem mem_bottom_track_35 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size8_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size8_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size8_25_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size8_25_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size5 mux_top_track_36 (
		.in({chanx_right_in[22], chanx_right_in[43], chany_bottom_in[43], chanx_left_in[30], chanx_left_in[43]}),
		.sram(mux_tree_tapbuf_L1SB_size5_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size5_0_sram_inv[0:2]),
		.out(chany_top_out[18]));

	mux_tree_tapbuf_L1SB_size5 mux_bottom_track_37 (
		.in({chany_top_in[43], chanx_right_in[22], chanx_right_in[43], chanx_left_in[22], chanx_left_in[43]}),
		.sram(mux_tree_tapbuf_L1SB_size5_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size5_1_sram_inv[0:2]),
		.out(chany_bottom_out[18]));

	mux_tree_tapbuf_L1SB_size5_mem mem_top_track_36 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size8_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size5_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size5_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size5_0_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size5_mem mem_bottom_track_37 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size8_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size5_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size5_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size5_1_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size5 mux_top_track_38 (
		.in({chanx_right_in[26], chanx_right_in[44], chany_bottom_in[44], chanx_left_in[26], chanx_left_in[44]}),
		.sram(mux_tree_tapbuf_L4SB_size5_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_0_sram_inv[0:2]),
		.out(chany_top_out[19]));

	mux_tree_tapbuf_L4SB_size5 mux_top_track_46 (
		.in({chanx_right_in[30], chanx_right_in[45], chany_bottom_in[45], chanx_left_in[22], chanx_left_in[45]}),
		.sram(mux_tree_tapbuf_L4SB_size5_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_1_sram_inv[0:2]),
		.out(chany_top_out[23]));

	mux_tree_tapbuf_L4SB_size5 mux_top_track_54 (
		.in({chanx_right_in[34], chanx_right_in[47], chany_bottom_in[47], chanx_left_in[18], chanx_left_in[47]}),
		.sram(mux_tree_tapbuf_L4SB_size5_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_2_sram_inv[0:2]),
		.out(chany_top_out[27]));

	mux_tree_tapbuf_L4SB_size5 mux_top_track_62 (
		.in({chanx_right_in[38], chanx_right_in[48], chany_bottom_in[48], chanx_left_in[17], chanx_left_in[48]}),
		.sram(mux_tree_tapbuf_L4SB_size5_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_3_sram_inv[0:2]),
		.out(chany_top_out[31]));

	mux_tree_tapbuf_L4SB_size5 mux_top_track_70 (
		.in({chanx_right_in[42], chanx_right_in[49], chany_bottom_in[49], chanx_left_in[16], chanx_left_in[49]}),
		.sram(mux_tree_tapbuf_L4SB_size5_4_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_4_sram_inv[0:2]),
		.out(chany_top_out[35]));

	mux_tree_tapbuf_L4SB_size5 mux_top_track_78 (
		.in({chanx_right_in[46], chanx_right_in[51], chany_bottom_in[51], chanx_left_in[15], chanx_left_in[51]}),
		.sram(mux_tree_tapbuf_L4SB_size5_5_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_5_sram_inv[0:2]),
		.out(chany_top_out[39]));

	mux_tree_tapbuf_L4SB_size5 mux_top_track_86 (
		.in({chanx_right_in[50], chanx_right_in[52], chany_bottom_in[52], chanx_left_in[14], chanx_left_in[52]}),
		.sram(mux_tree_tapbuf_L4SB_size5_6_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_6_sram_inv[0:2]),
		.out(chany_top_out[43]));

	mux_tree_tapbuf_L4SB_size5 mux_top_track_94 (
		.in({chanx_right_in[53:54], chany_bottom_in[53], chanx_left_in[13], chanx_left_in[53]}),
		.sram(mux_tree_tapbuf_L4SB_size5_7_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_7_sram_inv[0:2]),
		.out(chany_top_out[47]));

	mux_tree_tapbuf_L4SB_size5 mux_top_track_102 (
		.in({chanx_right_in[55], chanx_right_in[58], chany_bottom_in[55], chanx_left_in[12], chanx_left_in[55]}),
		.sram(mux_tree_tapbuf_L4SB_size5_8_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_8_sram_inv[0:2]),
		.out(chany_top_out[51]));

	mux_tree_tapbuf_L4SB_size5 mux_top_track_110 (
		.in({chanx_right_in[56], chanx_right_in[62], chany_bottom_in[56], chanx_left_in[11], chanx_left_in[56]}),
		.sram(mux_tree_tapbuf_L4SB_size5_9_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_9_sram_inv[0:2]),
		.out(chany_top_out[55]));

	mux_tree_tapbuf_L4SB_size5 mux_top_track_118 (
		.in({chanx_right_in[57], chanx_right_in[66], chany_bottom_in[57], chanx_left_in[10], chanx_left_in[57]}),
		.sram(mux_tree_tapbuf_L4SB_size5_10_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_10_sram_inv[0:2]),
		.out(chany_top_out[59]));

	mux_tree_tapbuf_L4SB_size5 mux_top_track_126 (
		.in({chanx_right_in[59], chanx_right_in[70], chany_bottom_in[59], chanx_left_in[9], chanx_left_in[59]}),
		.sram(mux_tree_tapbuf_L4SB_size5_11_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_11_sram_inv[0:2]),
		.out(chany_top_out[63]));

	mux_tree_tapbuf_L4SB_size5 mux_top_track_134 (
		.in({chanx_right_in[60], chanx_right_in[74], chany_bottom_in[60], chanx_left_in[8], chanx_left_in[60]}),
		.sram(mux_tree_tapbuf_L4SB_size5_12_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_12_sram_inv[0:2]),
		.out(chany_top_out[67]));

	mux_tree_tapbuf_L4SB_size5 mux_top_track_142 (
		.in({chanx_right_in[61], chanx_right_in[78], chany_bottom_in[61], chanx_left_in[7], chanx_left_in[61]}),
		.sram(mux_tree_tapbuf_L4SB_size5_13_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_13_sram_inv[0:2]),
		.out(chany_top_out[71]));

	mux_tree_tapbuf_L4SB_size5 mux_top_track_150 (
		.in({chanx_right_in[63], chanx_right_in[82], chany_bottom_in[63], chanx_left_in[6], chanx_left_in[63]}),
		.sram(mux_tree_tapbuf_L4SB_size5_14_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_14_sram_inv[0:2]),
		.out(chany_top_out[75]));

	mux_tree_tapbuf_L4SB_size5 mux_top_track_158 (
		.in({chanx_right_in[64], chanx_right_in[86], chany_bottom_in[64], chanx_left_in[5], chanx_left_in[64]}),
		.sram(mux_tree_tapbuf_L4SB_size5_15_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_15_sram_inv[0:2]),
		.out(chany_top_out[79]));

	mux_tree_tapbuf_L4SB_size5 mux_top_track_166 (
		.in({chanx_right_in[65], chanx_right_in[90], chany_bottom_in[65], chanx_left_in[4], chanx_left_in[65]}),
		.sram(mux_tree_tapbuf_L4SB_size5_16_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_16_sram_inv[0:2]),
		.out(chany_top_out[83]));

	mux_tree_tapbuf_L4SB_size5 mux_top_track_174 (
		.in({chanx_right_in[67], chanx_right_in[94], chany_bottom_in[67], chanx_left_in[3], chanx_left_in[67]}),
		.sram(mux_tree_tapbuf_L4SB_size5_17_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_17_sram_inv[0:2]),
		.out(chany_top_out[87]));

	mux_tree_tapbuf_L4SB_size5 mux_top_track_182 (
		.in({chanx_right_in[68], chanx_right_in[95], chany_bottom_in[68], chanx_left_in[2], chanx_left_in[68]}),
		.sram(mux_tree_tapbuf_L4SB_size5_18_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_18_sram_inv[0:2]),
		.out(chany_top_out[91]));

	mux_tree_tapbuf_L4SB_size5 mux_top_track_190 (
		.in({chanx_right_in[0], chanx_right_in[69], chany_bottom_in[69], chanx_left_in[1], chanx_left_in[69]}),
		.sram(mux_tree_tapbuf_L4SB_size5_19_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_19_sram_inv[0:2]),
		.out(chany_top_out[95]));

	mux_tree_tapbuf_L4SB_size5_mem mem_top_track_38 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size5_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size5_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size5_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_0_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size5_mem mem_top_track_46 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size5_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size5_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size5_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_1_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size5_mem mem_top_track_54 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size5_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size5_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size5_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_2_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size5_mem mem_top_track_62 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size5_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size5_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size5_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_3_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size5_mem mem_top_track_70 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size5_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size5_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size5_4_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_4_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size5_mem mem_top_track_78 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size5_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size5_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size5_5_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_5_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size5_mem mem_top_track_86 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size5_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size5_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size5_6_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_6_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size5_mem mem_top_track_94 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size5_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size5_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size5_7_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_7_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size5_mem mem_top_track_102 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size5_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size5_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size5_8_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_8_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size5_mem mem_top_track_110 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size5_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size5_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size5_9_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_9_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size5_mem mem_top_track_118 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size5_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size5_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size5_10_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_10_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size5_mem mem_top_track_126 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size5_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size5_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size5_11_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_11_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size5_mem mem_top_track_134 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size5_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size5_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size5_12_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_12_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size5_mem mem_top_track_142 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size5_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size5_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size5_13_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_13_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size5_mem mem_top_track_150 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size5_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size5_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size5_14_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_14_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size5_mem mem_top_track_158 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size5_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size5_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size5_15_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_15_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size5_mem mem_top_track_166 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size5_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size5_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size5_16_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_16_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size5_mem mem_top_track_174 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size5_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size5_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size5_17_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_17_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size5_mem mem_top_track_182 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size5_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size5_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size5_18_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_18_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size5_mem mem_top_track_190 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size5_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size5_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size5_19_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_19_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size10 mux_right_track_0 (
		.in({chany_top_in[19], chany_top_in[71], chany_top_in[95], right_top_grid_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_19__pin_a2f_o_0_, chany_bottom_in[19], chany_bottom_in[71], chany_bottom_in[94], chanx_left_in[19], chanx_left_in[71]}),
		.sram(mux_tree_tapbuf_L1SB_size10_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size10_0_sram_inv[0:3]),
		.out(chanx_right_out[0]));

	mux_tree_tapbuf_L1SB_size10 mux_left_track_1 (
		.in({chany_top_in[0], chany_top_in[19], chany_top_in[71], chanx_right_in[19], chanx_right_in[71], chany_bottom_in[19], chany_bottom_in[71], chany_bottom_in[95], left_top_grid_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_19__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L1SB_size10_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size10_1_sram_inv[0:3]),
		.out(chanx_left_out[0]));

	mux_tree_tapbuf_L1SB_size10 mux_left_track_3 (
		.in({chany_top_in[20], chany_top_in[72], chany_top_in[95], chanx_right_in[20], chanx_right_in[72], chany_bottom_in[0], chany_bottom_in[20], chany_bottom_in[72], left_top_grid_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_}),
		.sram(mux_tree_tapbuf_L1SB_size10_2_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size10_2_sram_inv[0:3]),
		.out(chanx_left_out[1]));

	mux_tree_tapbuf_L1SB_size10 mux_left_track_5 (
		.in({chany_top_in[21], chany_top_in[73], chany_top_in[94], chanx_right_in[21], chanx_right_in[73], chany_bottom_in[1], chany_bottom_in[21], chany_bottom_in[73], left_top_grid_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_}),
		.sram(mux_tree_tapbuf_L1SB_size10_3_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size10_3_sram_inv[0:3]),
		.out(chanx_left_out[2]));

	mux_tree_tapbuf_L1SB_size10 mux_left_track_7 (
		.in({chany_top_in[23], chany_top_in[75], chany_top_in[90], chanx_right_in[23], chanx_right_in[75], chany_bottom_in[2], chany_bottom_in[23], chany_bottom_in[75], left_top_grid_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_L1SB_size10_4_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size10_4_sram_inv[0:3]),
		.out(chanx_left_out[3]));

	mux_tree_tapbuf_L1SB_size10 mux_left_track_9 (
		.in({chany_top_in[24], chany_top_in[76], chany_top_in[86], chanx_right_in[24], chanx_right_in[76], chany_bottom_in[3], chany_bottom_in[24], chany_bottom_in[76], left_top_grid_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_}),
		.sram(mux_tree_tapbuf_L1SB_size10_5_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size10_5_sram_inv[0:3]),
		.out(chanx_left_out[4]));

	mux_tree_tapbuf_L1SB_size10 mux_left_track_11 (
		.in({chany_top_in[25], chany_top_in[77], chany_top_in[82], chanx_right_in[25], chanx_right_in[77], chany_bottom_in[4], chany_bottom_in[25], chany_bottom_in[77], left_top_grid_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_}),
		.sram(mux_tree_tapbuf_L1SB_size10_6_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size10_6_sram_inv[0:3]),
		.out(chanx_left_out[5]));

	mux_tree_tapbuf_L1SB_size10 mux_left_track_13 (
		.in({chany_top_in[27], chany_top_in[78:79], chanx_right_in[27], chanx_right_in[79], chany_bottom_in[5], chany_bottom_in[27], chany_bottom_in[79], left_top_grid_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_}),
		.sram(mux_tree_tapbuf_L1SB_size10_7_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size10_7_sram_inv[0:3]),
		.out(chanx_left_out[6]));

	mux_tree_tapbuf_L1SB_size10 mux_left_track_15 (
		.in({chany_top_in[28], chany_top_in[74], chany_top_in[80], chanx_right_in[28], chanx_right_in[80], chany_bottom_in[6], chany_bottom_in[28], chany_bottom_in[80], left_top_grid_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_}),
		.sram(mux_tree_tapbuf_L1SB_size10_8_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size10_8_sram_inv[0:3]),
		.out(chanx_left_out[7]));

	mux_tree_tapbuf_L1SB_size10 mux_left_track_17 (
		.in({chany_top_in[29], chany_top_in[70], chany_top_in[81], chanx_right_in[29], chanx_right_in[81], chany_bottom_in[7], chany_bottom_in[29], chany_bottom_in[81], left_top_grid_bottom_width_0_height_0_subtile_8__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_}),
		.sram(mux_tree_tapbuf_L1SB_size10_9_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size10_9_sram_inv[0:3]),
		.out(chanx_left_out[8]));

	mux_tree_tapbuf_L1SB_size10 mux_left_track_19 (
		.in({chany_top_in[31], chany_top_in[66], chany_top_in[83], chanx_right_in[31], chanx_right_in[83], chany_bottom_in[8], chany_bottom_in[31], chany_bottom_in[83], left_top_grid_bottom_width_0_height_0_subtile_9__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_}),
		.sram(mux_tree_tapbuf_L1SB_size10_10_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size10_10_sram_inv[0:3]),
		.out(chanx_left_out[9]));

	mux_tree_tapbuf_L1SB_size10 mux_left_track_21 (
		.in({chany_top_in[32], chany_top_in[62], chany_top_in[84], chanx_right_in[32], chanx_right_in[84], chany_bottom_in[9], chany_bottom_in[32], chany_bottom_in[84], left_top_grid_bottom_width_0_height_0_subtile_10__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_}),
		.sram(mux_tree_tapbuf_L1SB_size10_11_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size10_11_sram_inv[0:3]),
		.out(chanx_left_out[10]));

	mux_tree_tapbuf_L1SB_size10_mem mem_right_track_0 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size5_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size10_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size10_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size10_0_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size10_mem mem_left_track_1 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size7_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size10_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size10_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size10_1_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size10_mem mem_left_track_3 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size10_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size10_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size10_2_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size10_2_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size10_mem mem_left_track_5 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size10_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size10_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size10_3_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size10_3_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size10_mem mem_left_track_7 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size10_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size10_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size10_4_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size10_4_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size10_mem mem_left_track_9 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size10_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size10_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size10_5_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size10_5_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size10_mem mem_left_track_11 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size10_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size10_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size10_6_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size10_6_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size10_mem mem_left_track_13 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size10_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size10_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size10_7_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size10_7_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size10_mem mem_left_track_15 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size10_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size10_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size10_8_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size10_8_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size10_mem mem_left_track_17 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size10_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size10_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size10_9_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size10_9_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size10_mem mem_left_track_19 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size10_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size10_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size10_10_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size10_10_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size10_mem mem_left_track_21 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size10_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size10_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size10_11_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size10_11_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9 mux_right_track_2 (
		.in({chany_top_in[0], chany_top_in[20], chany_top_in[72], right_top_grid_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_, chany_bottom_in[20], chany_bottom_in[72], chany_bottom_in[90], chanx_left_in[20], chanx_left_in[72]}),
		.sram(mux_tree_tapbuf_L1SB_size9_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_0_sram_inv[0:3]),
		.out(chanx_right_out[1]));

	mux_tree_tapbuf_L1SB_size9 mux_right_track_4 (
		.in({chany_top_in[1], chany_top_in[21], chany_top_in[73], right_top_grid_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_, chany_bottom_in[21], chany_bottom_in[73], chany_bottom_in[86], chanx_left_in[21], chanx_left_in[73]}),
		.sram(mux_tree_tapbuf_L1SB_size9_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_1_sram_inv[0:3]),
		.out(chanx_right_out[2]));

	mux_tree_tapbuf_L1SB_size9 mux_right_track_6 (
		.in({chany_top_in[2], chany_top_in[23], chany_top_in[75], right_top_grid_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_, chany_bottom_in[23], chany_bottom_in[75], chany_bottom_in[82], chanx_left_in[23], chanx_left_in[75]}),
		.sram(mux_tree_tapbuf_L1SB_size9_2_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_2_sram_inv[0:3]),
		.out(chanx_right_out[3]));

	mux_tree_tapbuf_L1SB_size9 mux_right_track_8 (
		.in({chany_top_in[3], chany_top_in[24], chany_top_in[76], right_top_grid_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_, chany_bottom_in[24], chany_bottom_in[76], chany_bottom_in[78], chanx_left_in[24], chanx_left_in[76]}),
		.sram(mux_tree_tapbuf_L1SB_size9_3_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_3_sram_inv[0:3]),
		.out(chanx_right_out[4]));

	mux_tree_tapbuf_L1SB_size9 mux_right_track_10 (
		.in({chany_top_in[4], chany_top_in[25], chany_top_in[77], right_top_grid_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_, chany_bottom_in[25], chany_bottom_in[74], chany_bottom_in[77], chanx_left_in[25], chanx_left_in[77]}),
		.sram(mux_tree_tapbuf_L1SB_size9_4_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_4_sram_inv[0:3]),
		.out(chanx_right_out[5]));

	mux_tree_tapbuf_L1SB_size9 mux_right_track_12 (
		.in({chany_top_in[5], chany_top_in[27], chany_top_in[79], right_top_grid_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_, chany_bottom_in[27], chany_bottom_in[70], chany_bottom_in[79], chanx_left_in[27], chanx_left_in[79]}),
		.sram(mux_tree_tapbuf_L1SB_size9_5_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_5_sram_inv[0:3]),
		.out(chanx_right_out[6]));

	mux_tree_tapbuf_L1SB_size9 mux_right_track_14 (
		.in({chany_top_in[6], chany_top_in[28], chany_top_in[80], right_top_grid_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_, chany_bottom_in[28], chany_bottom_in[66], chany_bottom_in[80], chanx_left_in[28], chanx_left_in[80]}),
		.sram(mux_tree_tapbuf_L1SB_size9_6_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_6_sram_inv[0:3]),
		.out(chanx_right_out[7]));

	mux_tree_tapbuf_L1SB_size9 mux_right_track_16 (
		.in({chany_top_in[7], chany_top_in[29], chany_top_in[81], right_top_grid_bottom_width_0_height_0_subtile_8__pin_a2f_o_0_, chany_bottom_in[29], chany_bottom_in[62], chany_bottom_in[81], chanx_left_in[29], chanx_left_in[81]}),
		.sram(mux_tree_tapbuf_L1SB_size9_7_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_7_sram_inv[0:3]),
		.out(chanx_right_out[8]));

	mux_tree_tapbuf_L1SB_size9 mux_right_track_18 (
		.in({chany_top_in[8], chany_top_in[31], chany_top_in[83], right_top_grid_bottom_width_0_height_0_subtile_9__pin_a2f_o_0_, chany_bottom_in[31], chany_bottom_in[58], chany_bottom_in[83], chanx_left_in[31], chanx_left_in[83]}),
		.sram(mux_tree_tapbuf_L1SB_size9_8_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_8_sram_inv[0:3]),
		.out(chanx_right_out[9]));

	mux_tree_tapbuf_L1SB_size9 mux_right_track_20 (
		.in({chany_top_in[9], chany_top_in[32], chany_top_in[84], right_top_grid_bottom_width_0_height_0_subtile_10__pin_a2f_o_0_, chany_bottom_in[32], chany_bottom_in[54], chany_bottom_in[84], chanx_left_in[32], chanx_left_in[84]}),
		.sram(mux_tree_tapbuf_L1SB_size9_9_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_9_sram_inv[0:3]),
		.out(chanx_right_out[10]));

	mux_tree_tapbuf_L1SB_size9 mux_right_track_22 (
		.in({chany_top_in[10], chany_top_in[33], chany_top_in[85], right_top_grid_bottom_width_0_height_0_subtile_11__pin_a2f_o_0_, chany_bottom_in[33], chany_bottom_in[50], chany_bottom_in[85], chanx_left_in[33], chanx_left_in[85]}),
		.sram(mux_tree_tapbuf_L1SB_size9_10_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_10_sram_inv[0:3]),
		.out(chanx_right_out[11]));

	mux_tree_tapbuf_L1SB_size9 mux_right_track_24 (
		.in({chany_top_in[11], chany_top_in[35], chany_top_in[87], right_top_grid_bottom_width_0_height_0_subtile_12__pin_a2f_o_0_, chany_bottom_in[35], chany_bottom_in[46], chany_bottom_in[87], chanx_left_in[35], chanx_left_in[87]}),
		.sram(mux_tree_tapbuf_L1SB_size9_11_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_11_sram_inv[0:3]),
		.out(chanx_right_out[12]));

	mux_tree_tapbuf_L1SB_size9 mux_right_track_26 (
		.in({chany_top_in[12], chany_top_in[36], chany_top_in[88], right_top_grid_bottom_width_0_height_0_subtile_13__pin_a2f_o_0_, chany_bottom_in[36], chany_bottom_in[42], chany_bottom_in[88], chanx_left_in[36], chanx_left_in[88]}),
		.sram(mux_tree_tapbuf_L1SB_size9_12_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_12_sram_inv[0:3]),
		.out(chanx_right_out[13]));

	mux_tree_tapbuf_L1SB_size9 mux_right_track_28 (
		.in({chany_top_in[13], chany_top_in[37], chany_top_in[89], right_top_grid_bottom_width_0_height_0_subtile_14__pin_a2f_o_0_, chany_bottom_in[37:38], chany_bottom_in[89], chanx_left_in[37], chanx_left_in[89]}),
		.sram(mux_tree_tapbuf_L1SB_size9_13_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_13_sram_inv[0:3]),
		.out(chanx_right_out[14]));

	mux_tree_tapbuf_L1SB_size9 mux_right_track_30 (
		.in({chany_top_in[14], chany_top_in[39], chany_top_in[91], right_top_grid_bottom_width_0_height_0_subtile_15__pin_a2f_o_0_, chany_bottom_in[34], chany_bottom_in[39], chany_bottom_in[91], chanx_left_in[39], chanx_left_in[91]}),
		.sram(mux_tree_tapbuf_L1SB_size9_14_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_14_sram_inv[0:3]),
		.out(chanx_right_out[15]));

	mux_tree_tapbuf_L1SB_size9 mux_right_track_32 (
		.in({chany_top_in[15], chany_top_in[40], chany_top_in[92], right_top_grid_bottom_width_0_height_0_subtile_16__pin_a2f_o_0_, chany_bottom_in[30], chany_bottom_in[40], chany_bottom_in[92], chanx_left_in[40], chanx_left_in[92]}),
		.sram(mux_tree_tapbuf_L1SB_size9_15_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_15_sram_inv[0:3]),
		.out(chanx_right_out[16]));

	mux_tree_tapbuf_L1SB_size9 mux_right_track_34 (
		.in({chany_top_in[16], chany_top_in[41], chany_top_in[93], right_top_grid_bottom_width_0_height_0_subtile_17__pin_a2f_o_0_, chany_bottom_in[26], chany_bottom_in[41], chany_bottom_in[93], chanx_left_in[41], chanx_left_in[93]}),
		.sram(mux_tree_tapbuf_L1SB_size9_16_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_16_sram_inv[0:3]),
		.out(chanx_right_out[17]));

	mux_tree_tapbuf_L1SB_size9 mux_bottom_track_1 (
		.in({chany_top_in[19], chany_top_in[71], chanx_right_in[19], chanx_right_in[71], chanx_right_in[94], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_, chanx_left_in[1], chanx_left_in[19], chanx_left_in[71]}),
		.sram(mux_tree_tapbuf_L1SB_size9_17_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_17_sram_inv[0:3]),
		.out(chany_bottom_out[0]));

	mux_tree_tapbuf_L1SB_size9 mux_bottom_track_3 (
		.in({chany_top_in[20], chany_top_in[72], chanx_right_in[20], chanx_right_in[72], chanx_right_in[90], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_, chanx_left_in[2], chanx_left_in[20], chanx_left_in[72]}),
		.sram(mux_tree_tapbuf_L1SB_size9_18_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_18_sram_inv[0:3]),
		.out(chany_bottom_out[1]));

	mux_tree_tapbuf_L1SB_size9 mux_bottom_track_5 (
		.in({chany_top_in[21], chany_top_in[73], chanx_right_in[21], chanx_right_in[73], chanx_right_in[86], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_, chanx_left_in[3], chanx_left_in[21], chanx_left_in[73]}),
		.sram(mux_tree_tapbuf_L1SB_size9_19_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_19_sram_inv[0:3]),
		.out(chany_bottom_out[2]));

	mux_tree_tapbuf_L1SB_size9 mux_bottom_track_7 (
		.in({chany_top_in[23], chany_top_in[75], chanx_right_in[23], chanx_right_in[75], chanx_right_in[82], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, chanx_left_in[4], chanx_left_in[23], chanx_left_in[75]}),
		.sram(mux_tree_tapbuf_L1SB_size9_20_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_20_sram_inv[0:3]),
		.out(chany_bottom_out[3]));

	mux_tree_tapbuf_L1SB_size9 mux_bottom_track_9 (
		.in({chany_top_in[24], chany_top_in[76], chanx_right_in[24], chanx_right_in[76], chanx_right_in[78], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_, chanx_left_in[5], chanx_left_in[24], chanx_left_in[76]}),
		.sram(mux_tree_tapbuf_L1SB_size9_21_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_21_sram_inv[0:3]),
		.out(chany_bottom_out[4]));

	mux_tree_tapbuf_L1SB_size9 mux_bottom_track_11 (
		.in({chany_top_in[25], chany_top_in[77], chanx_right_in[25], chanx_right_in[74], chanx_right_in[77], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_, chanx_left_in[6], chanx_left_in[25], chanx_left_in[77]}),
		.sram(mux_tree_tapbuf_L1SB_size9_22_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_22_sram_inv[0:3]),
		.out(chany_bottom_out[5]));

	mux_tree_tapbuf_L1SB_size9 mux_bottom_track_13 (
		.in({chany_top_in[27], chany_top_in[79], chanx_right_in[27], chanx_right_in[70], chanx_right_in[79], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_16_, chanx_left_in[7], chanx_left_in[27], chanx_left_in[79]}),
		.sram(mux_tree_tapbuf_L1SB_size9_23_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_23_sram_inv[0:3]),
		.out(chany_bottom_out[6]));

	mux_tree_tapbuf_L1SB_size9 mux_bottom_track_15 (
		.in({chany_top_in[28], chany_top_in[80], chanx_right_in[28], chanx_right_in[66], chanx_right_in[80], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, chanx_left_in[8], chanx_left_in[28], chanx_left_in[80]}),
		.sram(mux_tree_tapbuf_L1SB_size9_24_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_24_sram_inv[0:3]),
		.out(chany_bottom_out[7]));

	mux_tree_tapbuf_L1SB_size9 mux_bottom_track_17 (
		.in({chany_top_in[29], chany_top_in[81], chanx_right_in[29], chanx_right_in[62], chanx_right_in[81], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_18_, chanx_left_in[9], chanx_left_in[29], chanx_left_in[81]}),
		.sram(mux_tree_tapbuf_L1SB_size9_25_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_25_sram_inv[0:3]),
		.out(chany_bottom_out[8]));

	mux_tree_tapbuf_L1SB_size9 mux_bottom_track_19 (
		.in({chany_top_in[31], chany_top_in[83], chanx_right_in[31], chanx_right_in[58], chanx_right_in[83], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_19_, chanx_left_in[10], chanx_left_in[31], chanx_left_in[83]}),
		.sram(mux_tree_tapbuf_L1SB_size9_26_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_26_sram_inv[0:3]),
		.out(chany_bottom_out[9]));

	mux_tree_tapbuf_L1SB_size9 mux_left_track_23 (
		.in({chany_top_in[33], chany_top_in[58], chany_top_in[85], chanx_right_in[33], chanx_right_in[85], chany_bottom_in[10], chany_bottom_in[33], chany_bottom_in[85], left_top_grid_bottom_width_0_height_0_subtile_11__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L1SB_size9_27_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_27_sram_inv[0:3]),
		.out(chanx_left_out[11]));

	mux_tree_tapbuf_L1SB_size9 mux_left_track_25 (
		.in({chany_top_in[35], chany_top_in[54], chany_top_in[87], chanx_right_in[35], chanx_right_in[87], chany_bottom_in[11], chany_bottom_in[35], chany_bottom_in[87], left_top_grid_bottom_width_0_height_0_subtile_12__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L1SB_size9_28_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_28_sram_inv[0:3]),
		.out(chanx_left_out[12]));

	mux_tree_tapbuf_L1SB_size9 mux_left_track_27 (
		.in({chany_top_in[36], chany_top_in[50], chany_top_in[88], chanx_right_in[36], chanx_right_in[88], chany_bottom_in[12], chany_bottom_in[36], chany_bottom_in[88], left_top_grid_bottom_width_0_height_0_subtile_13__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L1SB_size9_29_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_29_sram_inv[0:3]),
		.out(chanx_left_out[13]));

	mux_tree_tapbuf_L1SB_size9 mux_left_track_29 (
		.in({chany_top_in[37], chany_top_in[46], chany_top_in[89], chanx_right_in[37], chanx_right_in[89], chany_bottom_in[13], chany_bottom_in[37], chany_bottom_in[89], left_top_grid_bottom_width_0_height_0_subtile_14__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L1SB_size9_30_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_30_sram_inv[0:3]),
		.out(chanx_left_out[14]));

	mux_tree_tapbuf_L1SB_size9 mux_left_track_31 (
		.in({chany_top_in[39], chany_top_in[42], chany_top_in[91], chanx_right_in[39], chanx_right_in[91], chany_bottom_in[14], chany_bottom_in[39], chany_bottom_in[91], left_top_grid_bottom_width_0_height_0_subtile_15__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L1SB_size9_31_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_31_sram_inv[0:3]),
		.out(chanx_left_out[15]));

	mux_tree_tapbuf_L1SB_size9 mux_left_track_33 (
		.in({chany_top_in[38], chany_top_in[40], chany_top_in[92], chanx_right_in[40], chanx_right_in[92], chany_bottom_in[15], chany_bottom_in[40], chany_bottom_in[92], left_top_grid_bottom_width_0_height_0_subtile_16__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L1SB_size9_32_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_32_sram_inv[0:3]),
		.out(chanx_left_out[16]));

	mux_tree_tapbuf_L1SB_size9 mux_left_track_35 (
		.in({chany_top_in[34], chany_top_in[41], chany_top_in[93], chanx_right_in[41], chanx_right_in[93], chany_bottom_in[16], chany_bottom_in[41], chany_bottom_in[93], left_top_grid_bottom_width_0_height_0_subtile_17__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L1SB_size9_33_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L1SB_size9_33_sram_inv[0:3]),
		.out(chanx_left_out[17]));

	mux_tree_tapbuf_L1SB_size9_mem mem_right_track_2 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size10_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size9_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size9_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_0_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_right_track_4 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size9_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size9_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size9_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_1_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_right_track_6 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size9_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size9_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size9_2_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_2_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_right_track_8 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size9_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size9_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size9_3_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_3_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_right_track_10 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size9_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size9_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size9_4_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_4_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_right_track_12 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size9_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size9_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size9_5_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_5_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_right_track_14 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size9_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size9_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size9_6_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_6_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_right_track_16 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size9_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size9_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size9_7_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_7_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_right_track_18 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size9_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size9_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size9_8_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_8_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_right_track_20 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size9_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size9_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size9_9_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_9_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_right_track_22 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size9_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size9_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size9_10_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_10_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_right_track_24 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size9_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size9_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size9_11_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_11_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_right_track_26 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size9_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size9_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size9_12_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_12_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_right_track_28 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size9_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size9_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size9_13_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_13_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_right_track_30 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size9_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size9_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size9_14_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_14_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_right_track_32 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size9_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size9_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size9_15_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_15_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_right_track_34 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size9_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size9_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size9_16_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_16_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_bottom_track_1 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size9_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size9_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size9_17_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_17_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_bottom_track_3 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size9_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size9_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size9_18_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_18_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_bottom_track_5 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size9_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size9_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size9_19_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_19_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_bottom_track_7 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size9_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size9_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size9_20_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_20_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_bottom_track_9 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size9_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size9_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size9_21_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_21_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_bottom_track_11 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size9_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size9_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size9_22_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_22_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_bottom_track_13 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size9_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size9_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size9_23_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_23_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_bottom_track_15 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size9_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size9_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size9_24_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_24_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_bottom_track_17 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size9_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size9_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size9_25_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_25_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_bottom_track_19 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size9_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size9_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size9_26_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_26_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_left_track_23 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size10_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size9_mem_27_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size9_27_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_27_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_left_track_25 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size9_mem_27_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size9_mem_28_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size9_28_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_28_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_left_track_27 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size9_mem_28_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size9_mem_29_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size9_29_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_29_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_left_track_29 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size9_mem_29_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size9_mem_30_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size9_30_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_30_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_left_track_31 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size9_mem_30_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size9_mem_31_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size9_31_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_31_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_left_track_33 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size9_mem_31_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size9_mem_32_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size9_32_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_32_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size9_mem mem_left_track_35 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size9_mem_32_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size9_mem_33_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size9_33_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L1SB_size9_33_sram_inv[0:3]));

	mux_tree_tapbuf_L1SB_size6 mux_right_track_36 (
		.in({chany_top_in[17], chany_top_in[43], right_top_grid_bottom_width_0_height_0_subtile_18__pin_a2f_o_0_, chany_bottom_in[22], chany_bottom_in[43], chanx_left_in[43]}),
		.sram(mux_tree_tapbuf_L1SB_size6_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size6_0_sram_inv[0:2]),
		.out(chanx_right_out[18]));

	mux_tree_tapbuf_L1SB_size6 mux_left_track_37 (
		.in({chany_top_in[30], chany_top_in[43], chanx_right_in[43], chany_bottom_in[17], chany_bottom_in[43], left_top_grid_bottom_width_0_height_0_subtile_18__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L1SB_size6_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L1SB_size6_1_sram_inv[0:2]),
		.out(chanx_left_out[18]));

	mux_tree_tapbuf_L1SB_size6_mem mem_right_track_36 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size9_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size6_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size6_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size6_0_sram_inv[0:2]));

	mux_tree_tapbuf_L1SB_size6_mem mem_left_track_37 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size9_mem_33_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L1SB_size6_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_L1SB_size6_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L1SB_size6_1_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size9 mux_right_track_38 (
		.in({chany_top_in[18], chany_top_in[44], right_top_grid_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_8__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_14__pin_a2f_o_0_, chany_bottom_in[18], chany_bottom_in[44], chanx_left_in[44]}),
		.sram(mux_tree_tapbuf_L4SB_size9_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_0_sram_inv[0:3]),
		.out(chanx_right_out[19]));

	mux_tree_tapbuf_L4SB_size9 mux_right_track_46 (
		.in({chany_top_in[22], chany_top_in[45], right_top_grid_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_9__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_15__pin_a2f_o_0_, chany_bottom_in[17], chany_bottom_in[45], chanx_left_in[45]}),
		.sram(mux_tree_tapbuf_L4SB_size9_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_1_sram_inv[0:3]),
		.out(chanx_right_out[23]));

	mux_tree_tapbuf_L4SB_size9 mux_right_track_54 (
		.in({chany_top_in[26], chany_top_in[47], right_top_grid_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_10__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_16__pin_a2f_o_0_, chany_bottom_in[16], chany_bottom_in[47], chanx_left_in[47]}),
		.sram(mux_tree_tapbuf_L4SB_size9_2_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_2_sram_inv[0:3]),
		.out(chanx_right_out[27]));

	mux_tree_tapbuf_L4SB_size9 mux_right_track_62 (
		.in({chany_top_in[30], chany_top_in[48], right_top_grid_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_11__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_17__pin_a2f_o_0_, chany_bottom_in[15], chany_bottom_in[48], chanx_left_in[48]}),
		.sram(mux_tree_tapbuf_L4SB_size9_3_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_3_sram_inv[0:3]),
		.out(chanx_right_out[31]));

	mux_tree_tapbuf_L4SB_size9 mux_right_track_70 (
		.in({chany_top_in[34], chany_top_in[49], right_top_grid_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_12__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_18__pin_a2f_o_0_, chany_bottom_in[14], chany_bottom_in[49], chanx_left_in[49]}),
		.sram(mux_tree_tapbuf_L4SB_size9_4_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_4_sram_inv[0:3]),
		.out(chanx_right_out[35]));

	mux_tree_tapbuf_L4SB_size9 mux_right_track_78 (
		.in({chany_top_in[38], chany_top_in[51], right_top_grid_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_13__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_19__pin_a2f_o_0_, chany_bottom_in[13], chany_bottom_in[51], chanx_left_in[51]}),
		.sram(mux_tree_tapbuf_L4SB_size9_5_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_5_sram_inv[0:3]),
		.out(chanx_right_out[39]));

	mux_tree_tapbuf_L4SB_size9 mux_right_track_86 (
		.in({chany_top_in[42], chany_top_in[52], right_top_grid_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_8__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_14__pin_a2f_o_0_, chany_bottom_in[12], chany_bottom_in[52], chanx_left_in[52]}),
		.sram(mux_tree_tapbuf_L4SB_size9_6_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_6_sram_inv[0:3]),
		.out(chanx_right_out[43]));

	mux_tree_tapbuf_L4SB_size9 mux_right_track_94 (
		.in({chany_top_in[46], chany_top_in[53], right_top_grid_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_9__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_15__pin_a2f_o_0_, chany_bottom_in[11], chany_bottom_in[53], chanx_left_in[53]}),
		.sram(mux_tree_tapbuf_L4SB_size9_7_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_7_sram_inv[0:3]),
		.out(chanx_right_out[47]));

	mux_tree_tapbuf_L4SB_size9 mux_right_track_102 (
		.in({chany_top_in[50], chany_top_in[55], right_top_grid_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_8__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_10__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_16__pin_a2f_o_0_, chany_bottom_in[10], chany_bottom_in[55], chanx_left_in[55]}),
		.sram(mux_tree_tapbuf_L4SB_size9_8_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_8_sram_inv[0:3]),
		.out(chanx_right_out[51]));

	mux_tree_tapbuf_L4SB_size9 mux_right_track_110 (
		.in({chany_top_in[54], chany_top_in[56], right_top_grid_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_9__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_11__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_17__pin_a2f_o_0_, chany_bottom_in[9], chany_bottom_in[56], chanx_left_in[56]}),
		.sram(mux_tree_tapbuf_L4SB_size9_9_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_9_sram_inv[0:3]),
		.out(chanx_right_out[55]));

	mux_tree_tapbuf_L4SB_size9 mux_right_track_118 (
		.in({chany_top_in[57:58], right_top_grid_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_10__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_12__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_18__pin_a2f_o_0_, chany_bottom_in[8], chany_bottom_in[57], chanx_left_in[57]}),
		.sram(mux_tree_tapbuf_L4SB_size9_10_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_10_sram_inv[0:3]),
		.out(chanx_right_out[59]));

	mux_tree_tapbuf_L4SB_size9 mux_right_track_126 (
		.in({chany_top_in[59], chany_top_in[62], right_top_grid_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_11__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_13__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_19__pin_a2f_o_0_, chany_bottom_in[7], chany_bottom_in[59], chanx_left_in[59]}),
		.sram(mux_tree_tapbuf_L4SB_size9_11_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_11_sram_inv[0:3]),
		.out(chanx_right_out[63]));

	mux_tree_tapbuf_L4SB_size9 mux_right_track_134 (
		.in({chany_top_in[60], chany_top_in[66], right_top_grid_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_12__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_14__pin_a2f_o_0_, chany_bottom_in[6], chany_bottom_in[60], chanx_left_in[60]}),
		.sram(mux_tree_tapbuf_L4SB_size9_12_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_12_sram_inv[0:3]),
		.out(chanx_right_out[67]));

	mux_tree_tapbuf_L4SB_size9 mux_right_track_142 (
		.in({chany_top_in[61], chany_top_in[70], right_top_grid_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_13__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_15__pin_a2f_o_0_, chany_bottom_in[5], chany_bottom_in[61], chanx_left_in[61]}),
		.sram(mux_tree_tapbuf_L4SB_size9_13_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_13_sram_inv[0:3]),
		.out(chanx_right_out[71]));

	mux_tree_tapbuf_L4SB_size9 mux_right_track_150 (
		.in({chany_top_in[63], chany_top_in[74], right_top_grid_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_8__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_14__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_16__pin_a2f_o_0_, chany_bottom_in[4], chany_bottom_in[63], chanx_left_in[63]}),
		.sram(mux_tree_tapbuf_L4SB_size9_14_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_14_sram_inv[0:3]),
		.out(chanx_right_out[75]));

	mux_tree_tapbuf_L4SB_size9 mux_right_track_158 (
		.in({chany_top_in[64], chany_top_in[78], right_top_grid_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_9__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_15__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_17__pin_a2f_o_0_, chany_bottom_in[3], chany_bottom_in[64], chanx_left_in[64]}),
		.sram(mux_tree_tapbuf_L4SB_size9_15_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_15_sram_inv[0:3]),
		.out(chanx_right_out[79]));

	mux_tree_tapbuf_L4SB_size9 mux_right_track_166 (
		.in({chany_top_in[65], chany_top_in[82], right_top_grid_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_10__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_16__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_18__pin_a2f_o_0_, chany_bottom_in[2], chany_bottom_in[65], chanx_left_in[65]}),
		.sram(mux_tree_tapbuf_L4SB_size9_16_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_16_sram_inv[0:3]),
		.out(chanx_right_out[83]));

	mux_tree_tapbuf_L4SB_size9 mux_right_track_174 (
		.in({chany_top_in[67], chany_top_in[86], right_top_grid_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_11__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_17__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_19__pin_a2f_o_0_, chany_bottom_in[1], chany_bottom_in[67], chanx_left_in[67]}),
		.sram(mux_tree_tapbuf_L4SB_size9_17_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_17_sram_inv[0:3]),
		.out(chanx_right_out[87]));

	mux_tree_tapbuf_L4SB_size9 mux_right_track_182 (
		.in({chany_top_in[68], chany_top_in[90], right_top_grid_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_12__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_18__pin_a2f_o_0_, chany_bottom_in[0], chany_bottom_in[68], chanx_left_in[68]}),
		.sram(mux_tree_tapbuf_L4SB_size9_18_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_18_sram_inv[0:3]),
		.out(chanx_right_out[91]));

	mux_tree_tapbuf_L4SB_size9 mux_right_track_190 (
		.in({chany_top_in[69], chany_top_in[94], right_top_grid_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_13__pin_a2f_o_0_, right_top_grid_bottom_width_0_height_0_subtile_19__pin_a2f_o_0_, chany_bottom_in[69], chany_bottom_in[95], chanx_left_in[69]}),
		.sram(mux_tree_tapbuf_L4SB_size9_19_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_19_sram_inv[0:3]),
		.out(chanx_right_out[95]));

	mux_tree_tapbuf_L4SB_size9_mem mem_right_track_38 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size6_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size9_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size9_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_0_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_right_track_46 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size9_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size9_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size9_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_1_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_right_track_54 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size9_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size9_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size9_2_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_2_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_right_track_62 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size9_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size9_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size9_3_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_3_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_right_track_70 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size9_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size9_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size9_4_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_4_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_right_track_78 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size9_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size9_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size9_5_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_5_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_right_track_86 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size9_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size9_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size9_6_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_6_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_right_track_94 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size9_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size9_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size9_7_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_7_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_right_track_102 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size9_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size9_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size9_8_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_8_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_right_track_110 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size9_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size9_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size9_9_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_9_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_right_track_118 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size9_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size9_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size9_10_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_10_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_right_track_126 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size9_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size9_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size9_11_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_11_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_right_track_134 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size9_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size9_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size9_12_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_12_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_right_track_142 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size9_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size9_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size9_13_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_13_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_right_track_150 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size9_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size9_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size9_14_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_14_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_right_track_158 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size9_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size9_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size9_15_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_15_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_right_track_166 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size9_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size9_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size9_16_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_16_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_right_track_174 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size9_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size9_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size9_17_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_17_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_right_track_182 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size9_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size9_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size9_18_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_18_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_right_track_190 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size9_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size9_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size9_19_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_19_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_39 (
		.in({chany_top_in[44], chanx_right_in[18], chanx_right_in[44], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_18_, chanx_left_in[26], chanx_left_in[44]}),
		.sram(mux_tree_tapbuf_L4SB_size8_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_0_sram_inv[0:2]),
		.out(chany_bottom_out[19]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_47 (
		.in({chany_top_in[45], chanx_right_in[17], chanx_right_in[45], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_19_, chanx_left_in[30], chanx_left_in[45]}),
		.sram(mux_tree_tapbuf_L4SB_size8_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_1_sram_inv[0:2]),
		.out(chany_bottom_out[23]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_87 (
		.in({chany_top_in[52], chanx_right_in[12], chanx_right_in[52], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_16_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_18_, chanx_left_in[50], chanx_left_in[52]}),
		.sram(mux_tree_tapbuf_L4SB_size8_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_2_sram_inv[0:2]),
		.out(chany_bottom_out[43]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_95 (
		.in({chany_top_in[53], chanx_right_in[11], chanx_right_in[53], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_19_, chanx_left_in[53:54]}),
		.sram(mux_tree_tapbuf_L4SB_size8_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_3_sram_inv[0:2]),
		.out(chany_bottom_out[47]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_39 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size5_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_0_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_47 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_1_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_87 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size7_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_2_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_95 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_3_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7 mux_bottom_track_55 (
		.in({chany_top_in[47], chanx_right_in[16], chanx_right_in[47], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_, chanx_left_in[34], chanx_left_in[47]}),
		.sram(mux_tree_tapbuf_L4SB_size7_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_0_sram_inv[0:2]),
		.out(chany_bottom_out[27]));

	mux_tree_tapbuf_L4SB_size7 mux_bottom_track_63 (
		.in({chany_top_in[48], chanx_right_in[15], chanx_right_in[48], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_, chanx_left_in[38], chanx_left_in[48]}),
		.sram(mux_tree_tapbuf_L4SB_size7_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_1_sram_inv[0:2]),
		.out(chany_bottom_out[31]));

	mux_tree_tapbuf_L4SB_size7 mux_bottom_track_71 (
		.in({chany_top_in[49], chanx_right_in[14], chanx_right_in[49], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_16_, chanx_left_in[42], chanx_left_in[49]}),
		.sram(mux_tree_tapbuf_L4SB_size7_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_2_sram_inv[0:2]),
		.out(chany_bottom_out[35]));

	mux_tree_tapbuf_L4SB_size7 mux_bottom_track_79 (
		.in({chany_top_in[51], chanx_right_in[13], chanx_right_in[51], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, chanx_left_in[46], chanx_left_in[51]}),
		.sram(mux_tree_tapbuf_L4SB_size7_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_3_sram_inv[0:2]),
		.out(chany_bottom_out[39]));

	mux_tree_tapbuf_L4SB_size7 mux_bottom_track_103 (
		.in({chany_top_in[55], chanx_right_in[10], chanx_right_in[55], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_18_, chanx_left_in[55], chanx_left_in[58]}),
		.sram(mux_tree_tapbuf_L4SB_size7_4_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_4_sram_inv[0:2]),
		.out(chany_bottom_out[51]));

	mux_tree_tapbuf_L4SB_size7 mux_bottom_track_111 (
		.in({chany_top_in[56], chanx_right_in[9], chanx_right_in[56], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_19_, chanx_left_in[56], chanx_left_in[62]}),
		.sram(mux_tree_tapbuf_L4SB_size7_5_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_5_sram_inv[0:2]),
		.out(chany_bottom_out[55]));

	mux_tree_tapbuf_L4SB_size7 mux_bottom_track_135 (
		.in({chany_top_in[60], chanx_right_in[6], chanx_right_in[60], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_16_, chanx_left_in[60], chanx_left_in[74]}),
		.sram(mux_tree_tapbuf_L4SB_size7_6_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_6_sram_inv[0:2]),
		.out(chany_bottom_out[67]));

	mux_tree_tapbuf_L4SB_size7 mux_bottom_track_143 (
		.in({chany_top_in[61], chanx_right_in[5], chanx_right_in[61], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, chanx_left_in[61], chanx_left_in[78]}),
		.sram(mux_tree_tapbuf_L4SB_size7_7_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_7_sram_inv[0:2]),
		.out(chany_bottom_out[71]));

	mux_tree_tapbuf_L4SB_size7 mux_bottom_track_151 (
		.in({chany_top_in[63], chanx_right_in[4], chanx_right_in[63], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_18_, chanx_left_in[63], chanx_left_in[82]}),
		.sram(mux_tree_tapbuf_L4SB_size7_8_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_8_sram_inv[0:2]),
		.out(chany_bottom_out[75]));

	mux_tree_tapbuf_L4SB_size7 mux_bottom_track_159 (
		.in({chany_top_in[64], chanx_right_in[3], chanx_right_in[64], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_19_, chanx_left_in[64], chanx_left_in[86]}),
		.sram(mux_tree_tapbuf_L4SB_size7_9_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_9_sram_inv[0:2]),
		.out(chany_bottom_out[79]));

	mux_tree_tapbuf_L4SB_size7 mux_bottom_track_183 (
		.in({chany_top_in[68], chanx_right_in[0], chanx_right_in[68], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_16_, chanx_left_in[68], chanx_left_in[95]}),
		.sram(mux_tree_tapbuf_L4SB_size7_10_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_10_sram_inv[0:2]),
		.out(chany_bottom_out[91]));

	mux_tree_tapbuf_L4SB_size7 mux_bottom_track_191 (
		.in({chany_top_in[69], chanx_right_in[69], chanx_right_in[95], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_, chanx_left_in[0], chanx_left_in[69]}),
		.sram(mux_tree_tapbuf_L4SB_size7_11_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_11_sram_inv[0:2]),
		.out(chany_bottom_out[95]));

	mux_tree_tapbuf_L4SB_size7_mem mem_bottom_track_55 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size7_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size7_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_0_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7_mem mem_bottom_track_63 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size7_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size7_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size7_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_1_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7_mem mem_bottom_track_71 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size7_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size7_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size7_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_2_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7_mem mem_bottom_track_79 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size7_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size7_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size7_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_3_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7_mem mem_bottom_track_103 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size7_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size7_4_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_4_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7_mem mem_bottom_track_111 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size7_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size7_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size7_5_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_5_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7_mem mem_bottom_track_135 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size6_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size7_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size7_6_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_6_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7_mem mem_bottom_track_143 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size7_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size7_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size7_7_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_7_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7_mem mem_bottom_track_151 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size7_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size7_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size7_8_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_8_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7_mem mem_bottom_track_159 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size7_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size7_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size7_9_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_9_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7_mem mem_bottom_track_183 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size6_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size7_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size7_10_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_10_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7_mem mem_bottom_track_191 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size7_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size7_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size7_11_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_11_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size6 mux_bottom_track_119 (
		.in({chany_top_in[57], chanx_right_in[8], chanx_right_in[57], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_, chanx_left_in[57], chanx_left_in[66]}),
		.sram(mux_tree_tapbuf_L4SB_size6_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size6_0_sram_inv[0:2]),
		.out(chany_bottom_out[59]));

	mux_tree_tapbuf_L4SB_size6 mux_bottom_track_127 (
		.in({chany_top_in[59], chanx_right_in[7], chanx_right_in[59], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_, chanx_left_in[59], chanx_left_in[70]}),
		.sram(mux_tree_tapbuf_L4SB_size6_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size6_1_sram_inv[0:2]),
		.out(chany_bottom_out[63]));

	mux_tree_tapbuf_L4SB_size6 mux_bottom_track_167 (
		.in({chany_top_in[65], chanx_right_in[2], chanx_right_in[65], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_, chanx_left_in[65], chanx_left_in[90]}),
		.sram(mux_tree_tapbuf_L4SB_size6_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size6_2_sram_inv[0:2]),
		.out(chany_bottom_out[83]));

	mux_tree_tapbuf_L4SB_size6 mux_bottom_track_175 (
		.in({chany_top_in[67], chanx_right_in[1], chanx_right_in[67], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_, chanx_left_in[67], chanx_left_in[94]}),
		.sram(mux_tree_tapbuf_L4SB_size6_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size6_3_sram_inv[0:2]),
		.out(chany_bottom_out[87]));

	mux_tree_tapbuf_L4SB_size6_mem mem_bottom_track_119 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size7_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size6_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size6_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size6_0_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size6_mem mem_bottom_track_127 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size6_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size6_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size6_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size6_1_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size6_mem mem_bottom_track_167 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size7_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size6_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size6_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size6_2_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size6_mem mem_bottom_track_175 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size6_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size6_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size6_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size6_3_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size12 mux_left_track_39 (
		.in({chany_top_in[26], chany_top_in[44], chanx_right_in[44], chany_bottom_in[18], chany_bottom_in[44], left_top_grid_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_8__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_14__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_}),
		.sram(mux_tree_tapbuf_L4SB_size12_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size12_0_sram_inv[0:3]),
		.out(chanx_left_out[19]));

	mux_tree_tapbuf_L4SB_size12 mux_left_track_47 (
		.in({chany_top_in[22], chany_top_in[45], chanx_right_in[45], chany_bottom_in[22], chany_bottom_in[45], left_top_grid_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_9__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_15__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_}),
		.sram(mux_tree_tapbuf_L4SB_size12_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size12_1_sram_inv[0:3]),
		.out(chanx_left_out[23]));

	mux_tree_tapbuf_L4SB_size12 mux_left_track_87 (
		.in({chany_top_in[14], chany_top_in[52], chanx_right_in[52], chany_bottom_in[42], chany_bottom_in[52], left_top_grid_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_8__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_14__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_}),
		.sram(mux_tree_tapbuf_L4SB_size12_2_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size12_2_sram_inv[0:3]),
		.out(chanx_left_out[43]));

	mux_tree_tapbuf_L4SB_size12 mux_left_track_95 (
		.in({chany_top_in[13], chany_top_in[53], chanx_right_in[53], chany_bottom_in[46], chany_bottom_in[53], left_top_grid_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_9__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_15__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_}),
		.sram(mux_tree_tapbuf_L4SB_size12_3_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size12_3_sram_inv[0:3]),
		.out(chanx_left_out[47]));

	mux_tree_tapbuf_L4SB_size12_mem mem_left_track_39 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L1SB_size6_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size12_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size12_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size12_0_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size12_mem mem_left_track_47 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size12_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size12_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size12_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size12_1_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size12_mem mem_left_track_87 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size11_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size12_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size12_2_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size12_2_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size12_mem mem_left_track_95 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size12_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size12_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size12_3_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size12_3_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size11 mux_left_track_55 (
		.in({chany_top_in[18], chany_top_in[47], chanx_right_in[47], chany_bottom_in[26], chany_bottom_in[47], left_top_grid_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_10__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_16__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_}),
		.sram(mux_tree_tapbuf_L4SB_size11_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size11_0_sram_inv[0:3]),
		.out(chanx_left_out[27]));

	mux_tree_tapbuf_L4SB_size11 mux_left_track_63 (
		.in({chany_top_in[17], chany_top_in[48], chanx_right_in[48], chany_bottom_in[30], chany_bottom_in[48], left_top_grid_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_11__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_17__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_}),
		.sram(mux_tree_tapbuf_L4SB_size11_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size11_1_sram_inv[0:3]),
		.out(chanx_left_out[31]));

	mux_tree_tapbuf_L4SB_size11 mux_left_track_71 (
		.in({chany_top_in[16], chany_top_in[49], chanx_right_in[49], chany_bottom_in[34], chany_bottom_in[49], left_top_grid_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_12__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_18__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_}),
		.sram(mux_tree_tapbuf_L4SB_size11_2_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size11_2_sram_inv[0:3]),
		.out(chanx_left_out[35]));

	mux_tree_tapbuf_L4SB_size11 mux_left_track_79 (
		.in({chany_top_in[15], chany_top_in[51], chanx_right_in[51], chany_bottom_in[38], chany_bottom_in[51], left_top_grid_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_13__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_19__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_}),
		.sram(mux_tree_tapbuf_L4SB_size11_3_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size11_3_sram_inv[0:3]),
		.out(chanx_left_out[39]));

	mux_tree_tapbuf_L4SB_size11 mux_left_track_103 (
		.in({chany_top_in[12], chany_top_in[55], chanx_right_in[55], chany_bottom_in[50], chany_bottom_in[55], left_top_grid_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_8__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_10__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_16__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_}),
		.sram(mux_tree_tapbuf_L4SB_size11_4_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size11_4_sram_inv[0:3]),
		.out(chanx_left_out[51]));

	mux_tree_tapbuf_L4SB_size11 mux_left_track_111 (
		.in({chany_top_in[11], chany_top_in[56], chanx_right_in[56], chany_bottom_in[54], chany_bottom_in[56], left_top_grid_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_9__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_11__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_17__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_}),
		.sram(mux_tree_tapbuf_L4SB_size11_5_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size11_5_sram_inv[0:3]),
		.out(chanx_left_out[55]));

	mux_tree_tapbuf_L4SB_size11 mux_left_track_135 (
		.in({chany_top_in[8], chany_top_in[60], chanx_right_in[60], chany_bottom_in[60], chany_bottom_in[66], left_top_grid_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_12__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_14__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_}),
		.sram(mux_tree_tapbuf_L4SB_size11_6_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size11_6_sram_inv[0:3]),
		.out(chanx_left_out[67]));

	mux_tree_tapbuf_L4SB_size11 mux_left_track_143 (
		.in({chany_top_in[7], chany_top_in[61], chanx_right_in[61], chany_bottom_in[61], chany_bottom_in[70], left_top_grid_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_13__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_15__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_}),
		.sram(mux_tree_tapbuf_L4SB_size11_7_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size11_7_sram_inv[0:3]),
		.out(chanx_left_out[71]));

	mux_tree_tapbuf_L4SB_size11 mux_left_track_151 (
		.in({chany_top_in[6], chany_top_in[63], chanx_right_in[63], chany_bottom_in[63], chany_bottom_in[74], left_top_grid_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_8__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_14__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_16__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_}),
		.sram(mux_tree_tapbuf_L4SB_size11_8_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size11_8_sram_inv[0:3]),
		.out(chanx_left_out[75]));

	mux_tree_tapbuf_L4SB_size11 mux_left_track_159 (
		.in({chany_top_in[5], chany_top_in[64], chanx_right_in[64], chany_bottom_in[64], chany_bottom_in[78], left_top_grid_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_9__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_15__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_17__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_}),
		.sram(mux_tree_tapbuf_L4SB_size11_9_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size11_9_sram_inv[0:3]),
		.out(chanx_left_out[79]));

	mux_tree_tapbuf_L4SB_size11 mux_left_track_183 (
		.in({chany_top_in[2], chany_top_in[68], chanx_right_in[68], chany_bottom_in[68], chany_bottom_in[90], left_top_grid_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_12__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_18__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_}),
		.sram(mux_tree_tapbuf_L4SB_size11_10_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size11_10_sram_inv[0:3]),
		.out(chanx_left_out[91]));

	mux_tree_tapbuf_L4SB_size11 mux_left_track_191 (
		.in({chany_top_in[1], chany_top_in[69], chanx_right_in[69], chany_bottom_in[69], chany_bottom_in[94], left_top_grid_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_13__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_19__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_}),
		.sram(mux_tree_tapbuf_L4SB_size11_11_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size11_11_sram_inv[0:3]),
		.out(chanx_left_out[95]));

	mux_tree_tapbuf_L4SB_size11_mem mem_left_track_55 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size12_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size11_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size11_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size11_0_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size11_mem mem_left_track_63 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size11_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size11_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size11_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size11_1_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size11_mem mem_left_track_71 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size11_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size11_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size11_2_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size11_2_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size11_mem mem_left_track_79 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size11_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size11_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size11_3_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size11_3_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size11_mem mem_left_track_103 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size12_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size11_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size11_4_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size11_4_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size11_mem mem_left_track_111 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size11_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size11_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size11_5_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size11_5_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size11_mem mem_left_track_135 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size10_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size11_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size11_6_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size11_6_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size11_mem mem_left_track_143 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size11_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size11_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size11_7_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size11_7_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size11_mem mem_left_track_151 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size11_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size11_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size11_8_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size11_8_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size11_mem mem_left_track_159 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size11_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size11_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size11_9_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size11_9_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size11_mem mem_left_track_183 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size10_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size11_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size11_10_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size11_10_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size11_mem mem_left_track_191 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size11_mem_10_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size11_11_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size11_11_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size10 mux_left_track_119 (
		.in({chany_top_in[10], chany_top_in[57], chanx_right_in[57], chany_bottom_in[57:58], left_top_grid_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_10__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_12__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_18__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_}),
		.sram(mux_tree_tapbuf_L4SB_size10_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size10_0_sram_inv[0:3]),
		.out(chanx_left_out[59]));

	mux_tree_tapbuf_L4SB_size10 mux_left_track_127 (
		.in({chany_top_in[9], chany_top_in[59], chanx_right_in[59], chany_bottom_in[59], chany_bottom_in[62], left_top_grid_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_11__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_13__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_19__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_}),
		.sram(mux_tree_tapbuf_L4SB_size10_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size10_1_sram_inv[0:3]),
		.out(chanx_left_out[63]));

	mux_tree_tapbuf_L4SB_size10 mux_left_track_167 (
		.in({chany_top_in[4], chany_top_in[65], chanx_right_in[65], chany_bottom_in[65], chany_bottom_in[82], left_top_grid_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_10__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_16__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_18__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_}),
		.sram(mux_tree_tapbuf_L4SB_size10_2_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size10_2_sram_inv[0:3]),
		.out(chanx_left_out[83]));

	mux_tree_tapbuf_L4SB_size10 mux_left_track_175 (
		.in({chany_top_in[3], chany_top_in[67], chanx_right_in[67], chany_bottom_in[67], chany_bottom_in[86], left_top_grid_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_11__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_17__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_19__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_}),
		.sram(mux_tree_tapbuf_L4SB_size10_3_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size10_3_sram_inv[0:3]),
		.out(chanx_left_out[87]));

	mux_tree_tapbuf_L4SB_size10_mem mem_left_track_119 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size11_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size10_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size10_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size10_0_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size10_mem mem_left_track_127 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size10_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size10_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size10_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size10_1_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size10_mem mem_left_track_167 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size11_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size10_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size10_2_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size10_2_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size10_mem mem_left_track_175 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size10_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size10_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size10_3_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size10_3_sram_inv[0:3]));

endmodule
// ----- END Verilog module for sb_3__7_ -----

//----- Default net type -----
`default_nettype none



