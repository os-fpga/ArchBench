//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Top-level Verilog module for FPGA
//	Author: Xifan TANG
//	Organization: University of Utah
//-------------------------------------------
//----- Time scale -----
`timescale 1ns / 1ps

//----- Default net type -----
`default_nettype wire

// ----- Verilog module for fpga_top -----
module fpga_top(clk,
                global_reset,
                scan_reset,
                test_en,
                scan_mode,
                scan_clk,
                config_enable,
                prog_clock,
                CFG_DONE,
                gfpga_pad_QL_PREIO_A2F,
                gfpga_pad_QL_PREIO_F2A,
                gfpga_pad_QL_PREIO_F2A_DEF0,
                gfpga_pad_QL_PREIO_F2A_DEF1,
                gfpga_pad_QL_PREIO_F2A_CLK,
                ccff_head,
                ccff_tail);
//----- GLOBAL PORTS -----
input [0:3] clk;
//----- GLOBAL PORTS -----
input [0:0] global_reset;
//----- GLOBAL PORTS -----
input [0:0] scan_reset;
//----- GLOBAL PORTS -----
input [0:0] test_en;
//----- GLOBAL PORTS -----
input [0:0] scan_mode;
//----- GLOBAL PORTS -----
input [0:0] scan_clk;
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_clock;
//----- GLOBAL PORTS -----
input [0:0] CFG_DONE;
//----- GPIN PORTS -----
input [0:639] gfpga_pad_QL_PREIO_A2F;
//----- GPOUT PORTS -----
output [0:639] gfpga_pad_QL_PREIO_F2A;
//----- GPOUT PORTS -----
output [0:639] gfpga_pad_QL_PREIO_F2A_DEF0;
//----- GPOUT PORTS -----
output [0:639] gfpga_pad_QL_PREIO_F2A_DEF1;
//----- GPOUT PORTS -----
output [0:639] gfpga_pad_QL_PREIO_F2A_CLK;
//----- INPUT PORTS -----
input [0:9] ccff_head;
//----- OUTPUT PORTS -----
output [0:9] ccff_tail;

//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:95] cbx_1__0__0_chanx_left_out;
wire [0:95] cbx_1__0__0_chanx_right_out;
wire [0:95] cbx_1__0__10_chanx_left_out;
wire [0:95] cbx_1__0__10_chanx_right_out;
wire [0:95] cbx_1__0__11_chanx_left_out;
wire [0:95] cbx_1__0__11_chanx_right_out;
wire [0:95] cbx_1__0__12_chanx_left_out;
wire [0:95] cbx_1__0__12_chanx_right_out;
wire [0:95] cbx_1__0__13_chanx_left_out;
wire [0:95] cbx_1__0__13_chanx_right_out;
wire [0:95] cbx_1__0__14_chanx_left_out;
wire [0:95] cbx_1__0__14_chanx_right_out;
wire [0:95] cbx_1__0__15_chanx_left_out;
wire [0:95] cbx_1__0__15_chanx_right_out;
wire [0:95] cbx_1__0__16_chanx_left_out;
wire [0:95] cbx_1__0__16_chanx_right_out;
wire [0:95] cbx_1__0__17_chanx_left_out;
wire [0:95] cbx_1__0__17_chanx_right_out;
wire [0:95] cbx_1__0__18_chanx_left_out;
wire [0:95] cbx_1__0__18_chanx_right_out;
wire [0:95] cbx_1__0__19_chanx_left_out;
wire [0:95] cbx_1__0__19_chanx_right_out;
wire [0:95] cbx_1__0__1_chanx_left_out;
wire [0:95] cbx_1__0__1_chanx_right_out;
wire [0:95] cbx_1__0__20_chanx_left_out;
wire [0:95] cbx_1__0__20_chanx_right_out;
wire [0:95] cbx_1__0__21_chanx_left_out;
wire [0:95] cbx_1__0__21_chanx_right_out;
wire [0:95] cbx_1__0__22_chanx_left_out;
wire [0:95] cbx_1__0__22_chanx_right_out;
wire [0:95] cbx_1__0__23_chanx_left_out;
wire [0:95] cbx_1__0__23_chanx_right_out;
wire [0:95] cbx_1__0__24_chanx_left_out;
wire [0:95] cbx_1__0__24_chanx_right_out;
wire [0:95] cbx_1__0__25_chanx_left_out;
wire [0:95] cbx_1__0__25_chanx_right_out;
wire [0:95] cbx_1__0__26_chanx_left_out;
wire [0:95] cbx_1__0__26_chanx_right_out;
wire [0:95] cbx_1__0__27_chanx_left_out;
wire [0:95] cbx_1__0__27_chanx_right_out;
wire [0:95] cbx_1__0__28_chanx_left_out;
wire [0:95] cbx_1__0__28_chanx_right_out;
wire [0:95] cbx_1__0__29_chanx_left_out;
wire [0:95] cbx_1__0__29_chanx_right_out;
wire [0:95] cbx_1__0__2_chanx_left_out;
wire [0:95] cbx_1__0__2_chanx_right_out;
wire [0:95] cbx_1__0__30_chanx_left_out;
wire [0:95] cbx_1__0__30_chanx_right_out;
wire [0:95] cbx_1__0__31_chanx_left_out;
wire [0:95] cbx_1__0__31_chanx_right_out;
wire [0:95] cbx_1__0__32_chanx_left_out;
wire [0:95] cbx_1__0__32_chanx_right_out;
wire [0:95] cbx_1__0__33_chanx_left_out;
wire [0:95] cbx_1__0__33_chanx_right_out;
wire [0:95] cbx_1__0__34_chanx_left_out;
wire [0:95] cbx_1__0__34_chanx_right_out;
wire [0:95] cbx_1__0__35_chanx_left_out;
wire [0:95] cbx_1__0__35_chanx_right_out;
wire [0:95] cbx_1__0__36_chanx_left_out;
wire [0:95] cbx_1__0__36_chanx_right_out;
wire [0:95] cbx_1__0__37_chanx_left_out;
wire [0:95] cbx_1__0__37_chanx_right_out;
wire [0:95] cbx_1__0__38_chanx_left_out;
wire [0:95] cbx_1__0__38_chanx_right_out;
wire [0:95] cbx_1__0__39_chanx_left_out;
wire [0:95] cbx_1__0__39_chanx_right_out;
wire [0:95] cbx_1__0__3_chanx_left_out;
wire [0:95] cbx_1__0__3_chanx_right_out;
wire [0:95] cbx_1__0__40_chanx_left_out;
wire [0:95] cbx_1__0__40_chanx_right_out;
wire [0:95] cbx_1__0__41_chanx_left_out;
wire [0:95] cbx_1__0__41_chanx_right_out;
wire [0:95] cbx_1__0__42_chanx_left_out;
wire [0:95] cbx_1__0__42_chanx_right_out;
wire [0:95] cbx_1__0__4_chanx_left_out;
wire [0:95] cbx_1__0__4_chanx_right_out;
wire [0:95] cbx_1__0__5_chanx_left_out;
wire [0:95] cbx_1__0__5_chanx_right_out;
wire [0:95] cbx_1__0__6_chanx_left_out;
wire [0:95] cbx_1__0__6_chanx_right_out;
wire [0:95] cbx_1__0__7_chanx_left_out;
wire [0:95] cbx_1__0__7_chanx_right_out;
wire [0:95] cbx_1__0__8_chanx_left_out;
wire [0:95] cbx_1__0__8_chanx_right_out;
wire [0:95] cbx_1__0__9_chanx_left_out;
wire [0:95] cbx_1__0__9_chanx_right_out;
wire [0:95] cbx_2__1__0_chanx_left_out;
wire [0:95] cbx_2__1__0_chanx_right_out;
wire [0:95] cbx_2__1__1_chanx_left_out;
wire [0:95] cbx_2__1__1_chanx_right_out;
wire [0:95] cbx_2__1__2_chanx_left_out;
wire [0:95] cbx_2__1__2_chanx_right_out;
wire [0:95] cbx_2__1__3_chanx_left_out;
wire [0:95] cbx_2__1__3_chanx_right_out;
wire [0:95] cbx_2__1__4_chanx_left_out;
wire [0:95] cbx_2__1__4_chanx_right_out;
wire [0:95] cbx_2__1__5_chanx_left_out;
wire [0:95] cbx_2__1__5_chanx_right_out;
wire [0:95] cbx_2__2__0_chanx_left_out;
wire [0:95] cbx_2__2__0_chanx_right_out;
wire [0:95] cbx_2__2__10_chanx_left_out;
wire [0:95] cbx_2__2__10_chanx_right_out;
wire [0:95] cbx_2__2__11_chanx_left_out;
wire [0:95] cbx_2__2__11_chanx_right_out;
wire [0:95] cbx_2__2__12_chanx_left_out;
wire [0:95] cbx_2__2__12_chanx_right_out;
wire [0:95] cbx_2__2__13_chanx_left_out;
wire [0:95] cbx_2__2__13_chanx_right_out;
wire [0:95] cbx_2__2__14_chanx_left_out;
wire [0:95] cbx_2__2__14_chanx_right_out;
wire [0:95] cbx_2__2__15_chanx_left_out;
wire [0:95] cbx_2__2__15_chanx_right_out;
wire [0:95] cbx_2__2__16_chanx_left_out;
wire [0:95] cbx_2__2__16_chanx_right_out;
wire [0:95] cbx_2__2__17_chanx_left_out;
wire [0:95] cbx_2__2__17_chanx_right_out;
wire [0:95] cbx_2__2__18_chanx_left_out;
wire [0:95] cbx_2__2__18_chanx_right_out;
wire [0:95] cbx_2__2__19_chanx_left_out;
wire [0:95] cbx_2__2__19_chanx_right_out;
wire [0:95] cbx_2__2__1_chanx_left_out;
wire [0:95] cbx_2__2__1_chanx_right_out;
wire [0:95] cbx_2__2__20_chanx_left_out;
wire [0:95] cbx_2__2__20_chanx_right_out;
wire [0:95] cbx_2__2__21_chanx_left_out;
wire [0:95] cbx_2__2__21_chanx_right_out;
wire [0:95] cbx_2__2__22_chanx_left_out;
wire [0:95] cbx_2__2__22_chanx_right_out;
wire [0:95] cbx_2__2__23_chanx_left_out;
wire [0:95] cbx_2__2__23_chanx_right_out;
wire [0:95] cbx_2__2__24_chanx_left_out;
wire [0:95] cbx_2__2__24_chanx_right_out;
wire [0:95] cbx_2__2__25_chanx_left_out;
wire [0:95] cbx_2__2__25_chanx_right_out;
wire [0:95] cbx_2__2__26_chanx_left_out;
wire [0:95] cbx_2__2__26_chanx_right_out;
wire [0:95] cbx_2__2__27_chanx_left_out;
wire [0:95] cbx_2__2__27_chanx_right_out;
wire [0:95] cbx_2__2__28_chanx_left_out;
wire [0:95] cbx_2__2__28_chanx_right_out;
wire [0:95] cbx_2__2__29_chanx_left_out;
wire [0:95] cbx_2__2__29_chanx_right_out;
wire [0:95] cbx_2__2__2_chanx_left_out;
wire [0:95] cbx_2__2__2_chanx_right_out;
wire [0:95] cbx_2__2__3_chanx_left_out;
wire [0:95] cbx_2__2__3_chanx_right_out;
wire [0:95] cbx_2__2__4_chanx_left_out;
wire [0:95] cbx_2__2__4_chanx_right_out;
wire [0:95] cbx_2__2__5_chanx_left_out;
wire [0:95] cbx_2__2__5_chanx_right_out;
wire [0:95] cbx_2__2__6_chanx_left_out;
wire [0:95] cbx_2__2__6_chanx_right_out;
wire [0:95] cbx_2__2__7_chanx_left_out;
wire [0:95] cbx_2__2__7_chanx_right_out;
wire [0:95] cbx_2__2__8_chanx_left_out;
wire [0:95] cbx_2__2__8_chanx_right_out;
wire [0:95] cbx_2__2__9_chanx_left_out;
wire [0:95] cbx_2__2__9_chanx_right_out;
wire [0:95] cbx_2__7__0_chanx_left_out;
wire [0:95] cbx_2__7__0_chanx_right_out;
wire [0:95] cbx_2__7__1_chanx_left_out;
wire [0:95] cbx_2__7__1_chanx_right_out;
wire [0:95] cbx_2__7__2_chanx_left_out;
wire [0:95] cbx_2__7__2_chanx_right_out;
wire [0:95] cbx_2__7__3_chanx_left_out;
wire [0:95] cbx_2__7__3_chanx_right_out;
wire [0:95] cbx_2__7__4_chanx_left_out;
wire [0:95] cbx_2__7__4_chanx_right_out;
wire [0:95] cbx_2__7__5_chanx_left_out;
wire [0:95] cbx_2__7__5_chanx_right_out;
wire [0:95] cbx_4__1__0_chanx_left_out;
wire [0:95] cbx_4__1__0_chanx_right_out;
wire [0:95] cbx_4__4__0_chanx_left_out;
wire [0:95] cbx_4__4__0_chanx_right_out;
wire [0:95] cbx_4__7__0_chanx_left_out;
wire [0:95] cbx_4__7__0_chanx_right_out;
wire [0:95] cbx_4__7__1_chanx_left_out;
wire [0:95] cbx_4__7__1_chanx_right_out;
wire [0:95] cbx_7__1__0_chanx_left_out;
wire [0:95] cbx_7__1__0_chanx_right_out;
wire [0:95] cby_0__1__0_chany_bottom_out;
wire [0:95] cby_0__1__0_chany_top_out;
wire [0:95] cby_0__1__10_chany_bottom_out;
wire [0:95] cby_0__1__10_chany_top_out;
wire [0:95] cby_0__1__11_chany_bottom_out;
wire [0:95] cby_0__1__11_chany_top_out;
wire [0:95] cby_0__1__12_chany_bottom_out;
wire [0:95] cby_0__1__12_chany_top_out;
wire [0:95] cby_0__1__13_chany_bottom_out;
wire [0:95] cby_0__1__13_chany_top_out;
wire [0:95] cby_0__1__14_chany_bottom_out;
wire [0:95] cby_0__1__14_chany_top_out;
wire [0:95] cby_0__1__15_chany_bottom_out;
wire [0:95] cby_0__1__15_chany_top_out;
wire [0:95] cby_0__1__16_chany_bottom_out;
wire [0:95] cby_0__1__16_chany_top_out;
wire [0:95] cby_0__1__17_chany_bottom_out;
wire [0:95] cby_0__1__17_chany_top_out;
wire [0:95] cby_0__1__18_chany_bottom_out;
wire [0:95] cby_0__1__18_chany_top_out;
wire [0:95] cby_0__1__19_chany_bottom_out;
wire [0:95] cby_0__1__19_chany_top_out;
wire [0:95] cby_0__1__1_chany_bottom_out;
wire [0:95] cby_0__1__1_chany_top_out;
wire [0:95] cby_0__1__20_chany_bottom_out;
wire [0:95] cby_0__1__20_chany_top_out;
wire [0:95] cby_0__1__21_chany_bottom_out;
wire [0:95] cby_0__1__21_chany_top_out;
wire [0:95] cby_0__1__22_chany_bottom_out;
wire [0:95] cby_0__1__22_chany_top_out;
wire [0:95] cby_0__1__23_chany_bottom_out;
wire [0:95] cby_0__1__23_chany_top_out;
wire [0:95] cby_0__1__24_chany_bottom_out;
wire [0:95] cby_0__1__24_chany_top_out;
wire [0:95] cby_0__1__25_chany_bottom_out;
wire [0:95] cby_0__1__25_chany_top_out;
wire [0:95] cby_0__1__26_chany_bottom_out;
wire [0:95] cby_0__1__26_chany_top_out;
wire [0:95] cby_0__1__27_chany_bottom_out;
wire [0:95] cby_0__1__27_chany_top_out;
wire [0:95] cby_0__1__28_chany_bottom_out;
wire [0:95] cby_0__1__28_chany_top_out;
wire [0:95] cby_0__1__29_chany_bottom_out;
wire [0:95] cby_0__1__29_chany_top_out;
wire [0:95] cby_0__1__2_chany_bottom_out;
wire [0:95] cby_0__1__2_chany_top_out;
wire [0:95] cby_0__1__3_chany_bottom_out;
wire [0:95] cby_0__1__3_chany_top_out;
wire [0:95] cby_0__1__4_chany_bottom_out;
wire [0:95] cby_0__1__4_chany_top_out;
wire [0:95] cby_0__1__5_chany_bottom_out;
wire [0:95] cby_0__1__5_chany_top_out;
wire [0:95] cby_0__1__6_chany_bottom_out;
wire [0:95] cby_0__1__6_chany_top_out;
wire [0:95] cby_0__1__7_chany_bottom_out;
wire [0:95] cby_0__1__7_chany_top_out;
wire [0:95] cby_0__1__8_chany_bottom_out;
wire [0:95] cby_0__1__8_chany_top_out;
wire [0:95] cby_0__1__9_chany_bottom_out;
wire [0:95] cby_0__1__9_chany_top_out;
wire [0:95] cby_1__1__0_chany_bottom_out;
wire [0:95] cby_1__1__0_chany_top_out;
wire [0:95] cby_1__1__1_chany_bottom_out;
wire [0:95] cby_1__1__1_chany_top_out;
wire [0:95] cby_1__1__2_chany_bottom_out;
wire [0:95] cby_1__1__2_chany_top_out;
wire [0:95] cby_1__1__3_chany_bottom_out;
wire [0:95] cby_1__1__3_chany_top_out;
wire [0:95] cby_1__1__4_chany_bottom_out;
wire [0:95] cby_1__1__4_chany_top_out;
wire [0:95] cby_1__1__5_chany_bottom_out;
wire [0:95] cby_1__1__5_chany_top_out;
wire [0:95] cby_1__1__6_chany_bottom_out;
wire [0:95] cby_1__1__6_chany_top_out;
wire [0:95] cby_1__1__7_chany_bottom_out;
wire [0:95] cby_1__1__7_chany_top_out;
wire [0:95] cby_2__2__0_chany_bottom_out;
wire [0:95] cby_2__2__0_chany_top_out;
wire [0:95] cby_2__2__10_chany_bottom_out;
wire [0:95] cby_2__2__10_chany_top_out;
wire [0:95] cby_2__2__11_chany_bottom_out;
wire [0:95] cby_2__2__11_chany_top_out;
wire [0:95] cby_2__2__12_chany_bottom_out;
wire [0:95] cby_2__2__12_chany_top_out;
wire [0:95] cby_2__2__13_chany_bottom_out;
wire [0:95] cby_2__2__13_chany_top_out;
wire [0:95] cby_2__2__14_chany_bottom_out;
wire [0:95] cby_2__2__14_chany_top_out;
wire [0:95] cby_2__2__15_chany_bottom_out;
wire [0:95] cby_2__2__15_chany_top_out;
wire [0:95] cby_2__2__16_chany_bottom_out;
wire [0:95] cby_2__2__16_chany_top_out;
wire [0:95] cby_2__2__17_chany_bottom_out;
wire [0:95] cby_2__2__17_chany_top_out;
wire [0:95] cby_2__2__18_chany_bottom_out;
wire [0:95] cby_2__2__18_chany_top_out;
wire [0:95] cby_2__2__19_chany_bottom_out;
wire [0:95] cby_2__2__19_chany_top_out;
wire [0:95] cby_2__2__1_chany_bottom_out;
wire [0:95] cby_2__2__1_chany_top_out;
wire [0:95] cby_2__2__20_chany_bottom_out;
wire [0:95] cby_2__2__20_chany_top_out;
wire [0:95] cby_2__2__21_chany_bottom_out;
wire [0:95] cby_2__2__21_chany_top_out;
wire [0:95] cby_2__2__22_chany_bottom_out;
wire [0:95] cby_2__2__22_chany_top_out;
wire [0:95] cby_2__2__23_chany_bottom_out;
wire [0:95] cby_2__2__23_chany_top_out;
wire [0:95] cby_2__2__24_chany_bottom_out;
wire [0:95] cby_2__2__24_chany_top_out;
wire [0:95] cby_2__2__25_chany_bottom_out;
wire [0:95] cby_2__2__25_chany_top_out;
wire [0:95] cby_2__2__26_chany_bottom_out;
wire [0:95] cby_2__2__26_chany_top_out;
wire [0:95] cby_2__2__27_chany_bottom_out;
wire [0:95] cby_2__2__27_chany_top_out;
wire [0:95] cby_2__2__28_chany_bottom_out;
wire [0:95] cby_2__2__28_chany_top_out;
wire [0:95] cby_2__2__29_chany_bottom_out;
wire [0:95] cby_2__2__29_chany_top_out;
wire [0:95] cby_2__2__2_chany_bottom_out;
wire [0:95] cby_2__2__2_chany_top_out;
wire [0:95] cby_2__2__3_chany_bottom_out;
wire [0:95] cby_2__2__3_chany_top_out;
wire [0:95] cby_2__2__4_chany_bottom_out;
wire [0:95] cby_2__2__4_chany_top_out;
wire [0:95] cby_2__2__5_chany_bottom_out;
wire [0:95] cby_2__2__5_chany_top_out;
wire [0:95] cby_2__2__6_chany_bottom_out;
wire [0:95] cby_2__2__6_chany_top_out;
wire [0:95] cby_2__2__7_chany_bottom_out;
wire [0:95] cby_2__2__7_chany_top_out;
wire [0:95] cby_2__2__8_chany_bottom_out;
wire [0:95] cby_2__2__8_chany_top_out;
wire [0:95] cby_2__2__9_chany_bottom_out;
wire [0:95] cby_2__2__9_chany_top_out;
wire [0:95] cby_4__2__0_chany_bottom_out;
wire [0:95] cby_4__2__0_chany_top_out;
wire [0:95] cby_4__2__1_chany_bottom_out;
wire [0:95] cby_4__2__1_chany_top_out;
wire [0:95] cby_4__3__0_chany_bottom_out;
wire [0:95] cby_4__3__0_chany_top_out;
wire [0:95] cby_4__3__1_chany_bottom_out;
wire [0:95] cby_4__3__1_chany_top_out;
wire [0:95] cby_4__4__0_chany_bottom_out;
wire [0:95] cby_4__4__0_chany_top_out;
wire [0:95] cby_4__4__1_chany_bottom_out;
wire [0:95] cby_4__4__1_chany_top_out;
wire [0:95] cby_7__2__0_chany_bottom_out;
wire [0:95] cby_7__2__0_chany_top_out;
wire [0:95] cby_7__3__0_chany_bottom_out;
wire [0:95] cby_7__3__0_chany_top_out;
wire [0:95] cby_7__4__0_chany_bottom_out;
wire [0:95] cby_7__4__0_chany_top_out;
wire [0:95] cby_7__5__0_chany_bottom_out;
wire [0:95] cby_7__5__0_chany_top_out;
wire [0:95] cby_7__6__0_chany_bottom_out;
wire [0:95] cby_7__6__0_chany_top_out;
wire [0:95] cby_7__7__0_chany_bottom_out;
wire [0:95] cby_7__7__0_chany_top_out;
wire [0:95] cby_9__1__0_chany_bottom_out;
wire [0:95] cby_9__1__0_chany_top_out;
wire [0:95] cby_9__1__1_chany_bottom_out;
wire [0:95] cby_9__1__1_chany_top_out;
wire [0:95] cby_9__2__0_chany_bottom_out;
wire [0:95] cby_9__2__0_chany_top_out;
wire [0:95] cby_9__2__1_chany_bottom_out;
wire [0:95] cby_9__2__1_chany_top_out;
wire [0:95] cby_9__2__2_chany_bottom_out;
wire [0:95] cby_9__2__2_chany_top_out;
wire [0:95] cby_9__2__3_chany_bottom_out;
wire [0:95] cby_9__2__3_chany_top_out;
wire [0:95] cby_9__2__4_chany_bottom_out;
wire [0:95] cby_9__2__4_chany_top_out;
wire [0:95] cby_9__2__5_chany_bottom_out;
wire [0:95] cby_9__2__5_chany_top_out;
wire [0:95] sb_0__0__0_chanx_right_out;
wire [0:95] sb_0__0__0_chany_top_out;
wire [0:95] sb_0__1__0_chanx_right_out;
wire [0:95] sb_0__1__0_chany_bottom_out;
wire [0:95] sb_0__1__0_chany_top_out;
wire [0:95] sb_0__1__1_chanx_right_out;
wire [0:95] sb_0__1__1_chany_bottom_out;
wire [0:95] sb_0__1__1_chany_top_out;
wire [0:95] sb_0__1__2_chanx_right_out;
wire [0:95] sb_0__1__2_chany_bottom_out;
wire [0:95] sb_0__1__2_chany_top_out;
wire [0:95] sb_0__1__3_chanx_right_out;
wire [0:95] sb_0__1__3_chany_bottom_out;
wire [0:95] sb_0__1__3_chany_top_out;
wire [0:95] sb_0__1__4_chanx_right_out;
wire [0:95] sb_0__1__4_chany_bottom_out;
wire [0:95] sb_0__1__4_chany_top_out;
wire [0:95] sb_0__1__5_chanx_right_out;
wire [0:95] sb_0__1__5_chany_bottom_out;
wire [0:95] sb_0__1__5_chany_top_out;
wire [0:95] sb_0__1__6_chanx_right_out;
wire [0:95] sb_0__1__6_chany_bottom_out;
wire [0:95] sb_0__1__6_chany_top_out;
wire [0:95] sb_0__8__0_chanx_right_out;
wire [0:95] sb_0__8__0_chany_bottom_out;
wire [0:95] sb_10__0__0_chanx_left_out;
wire [0:95] sb_10__0__0_chany_top_out;
wire [0:95] sb_10__1__0_chanx_left_out;
wire [0:95] sb_10__1__0_chany_bottom_out;
wire [0:95] sb_10__1__0_chany_top_out;
wire [0:95] sb_10__1__1_chanx_left_out;
wire [0:95] sb_10__1__1_chany_bottom_out;
wire [0:95] sb_10__1__1_chany_top_out;
wire [0:95] sb_10__1__2_chanx_left_out;
wire [0:95] sb_10__1__2_chany_bottom_out;
wire [0:95] sb_10__1__2_chany_top_out;
wire [0:95] sb_10__1__3_chanx_left_out;
wire [0:95] sb_10__1__3_chany_bottom_out;
wire [0:95] sb_10__1__3_chany_top_out;
wire [0:95] sb_10__1__4_chanx_left_out;
wire [0:95] sb_10__1__4_chany_bottom_out;
wire [0:95] sb_10__1__4_chany_top_out;
wire [0:95] sb_10__1__5_chanx_left_out;
wire [0:95] sb_10__1__5_chany_bottom_out;
wire [0:95] sb_10__1__5_chany_top_out;
wire [0:95] sb_10__1__6_chanx_left_out;
wire [0:95] sb_10__1__6_chany_bottom_out;
wire [0:95] sb_10__1__6_chany_top_out;
wire [0:95] sb_10__8__0_chanx_left_out;
wire [0:95] sb_10__8__0_chany_bottom_out;
wire [0:95] sb_1__0__0_chanx_left_out;
wire [0:95] sb_1__0__0_chanx_right_out;
wire [0:95] sb_1__0__0_chany_top_out;
wire [0:95] sb_1__0__1_chanx_left_out;
wire [0:95] sb_1__0__1_chanx_right_out;
wire [0:95] sb_1__0__1_chany_top_out;
wire [0:95] sb_1__1__0_chanx_left_out;
wire [0:95] sb_1__1__0_chanx_right_out;
wire [0:95] sb_1__1__0_chany_bottom_out;
wire [0:95] sb_1__1__0_chany_top_out;
wire [0:95] sb_1__2__0_chanx_left_out;
wire [0:95] sb_1__2__0_chanx_right_out;
wire [0:95] sb_1__2__0_chany_bottom_out;
wire [0:95] sb_1__2__0_chany_top_out;
wire [0:95] sb_1__2__1_chanx_left_out;
wire [0:95] sb_1__2__1_chanx_right_out;
wire [0:95] sb_1__2__1_chany_bottom_out;
wire [0:95] sb_1__2__1_chany_top_out;
wire [0:95] sb_1__2__2_chanx_left_out;
wire [0:95] sb_1__2__2_chanx_right_out;
wire [0:95] sb_1__2__2_chany_bottom_out;
wire [0:95] sb_1__2__2_chany_top_out;
wire [0:95] sb_1__2__3_chanx_left_out;
wire [0:95] sb_1__2__3_chanx_right_out;
wire [0:95] sb_1__2__3_chany_bottom_out;
wire [0:95] sb_1__2__3_chany_top_out;
wire [0:95] sb_1__2__4_chanx_left_out;
wire [0:95] sb_1__2__4_chanx_right_out;
wire [0:95] sb_1__2__4_chany_bottom_out;
wire [0:95] sb_1__2__4_chany_top_out;
wire [0:95] sb_1__7__0_chanx_left_out;
wire [0:95] sb_1__7__0_chanx_right_out;
wire [0:95] sb_1__7__0_chany_bottom_out;
wire [0:95] sb_1__7__0_chany_top_out;
wire [0:95] sb_1__8__0_chanx_left_out;
wire [0:95] sb_1__8__0_chanx_right_out;
wire [0:95] sb_1__8__0_chany_bottom_out;
wire [0:95] sb_1__8__1_chanx_left_out;
wire [0:95] sb_1__8__1_chanx_right_out;
wire [0:95] sb_1__8__1_chany_bottom_out;
wire [0:95] sb_2__0__0_chanx_left_out;
wire [0:95] sb_2__0__0_chanx_right_out;
wire [0:95] sb_2__0__0_chany_top_out;
wire [0:95] sb_2__0__1_chanx_left_out;
wire [0:95] sb_2__0__1_chanx_right_out;
wire [0:95] sb_2__0__1_chany_top_out;
wire [0:95] sb_2__0__2_chanx_left_out;
wire [0:95] sb_2__0__2_chanx_right_out;
wire [0:95] sb_2__0__2_chany_top_out;
wire [0:95] sb_2__0__3_chanx_left_out;
wire [0:95] sb_2__0__3_chanx_right_out;
wire [0:95] sb_2__0__3_chany_top_out;
wire [0:95] sb_2__0__4_chanx_left_out;
wire [0:95] sb_2__0__4_chanx_right_out;
wire [0:95] sb_2__0__4_chany_top_out;
wire [0:95] sb_2__0__5_chanx_left_out;
wire [0:95] sb_2__0__5_chanx_right_out;
wire [0:95] sb_2__0__5_chany_top_out;
wire [0:95] sb_2__0__6_chanx_left_out;
wire [0:95] sb_2__0__6_chanx_right_out;
wire [0:95] sb_2__0__6_chany_top_out;
wire [0:95] sb_2__1__0_chanx_left_out;
wire [0:95] sb_2__1__0_chanx_right_out;
wire [0:95] sb_2__1__0_chany_bottom_out;
wire [0:95] sb_2__1__0_chany_top_out;
wire [0:95] sb_2__1__1_chanx_left_out;
wire [0:95] sb_2__1__1_chanx_right_out;
wire [0:95] sb_2__1__1_chany_bottom_out;
wire [0:95] sb_2__1__1_chany_top_out;
wire [0:95] sb_2__1__2_chanx_left_out;
wire [0:95] sb_2__1__2_chanx_right_out;
wire [0:95] sb_2__1__2_chany_bottom_out;
wire [0:95] sb_2__1__2_chany_top_out;
wire [0:95] sb_2__1__3_chanx_left_out;
wire [0:95] sb_2__1__3_chanx_right_out;
wire [0:95] sb_2__1__3_chany_bottom_out;
wire [0:95] sb_2__1__3_chany_top_out;
wire [0:95] sb_2__2__0_chanx_left_out;
wire [0:95] sb_2__2__0_chanx_right_out;
wire [0:95] sb_2__2__0_chany_bottom_out;
wire [0:95] sb_2__2__0_chany_top_out;
wire [0:95] sb_2__2__10_chanx_left_out;
wire [0:95] sb_2__2__10_chanx_right_out;
wire [0:95] sb_2__2__10_chany_bottom_out;
wire [0:95] sb_2__2__10_chany_top_out;
wire [0:95] sb_2__2__11_chanx_left_out;
wire [0:95] sb_2__2__11_chanx_right_out;
wire [0:95] sb_2__2__11_chany_bottom_out;
wire [0:95] sb_2__2__11_chany_top_out;
wire [0:95] sb_2__2__12_chanx_left_out;
wire [0:95] sb_2__2__12_chanx_right_out;
wire [0:95] sb_2__2__12_chany_bottom_out;
wire [0:95] sb_2__2__12_chany_top_out;
wire [0:95] sb_2__2__13_chanx_left_out;
wire [0:95] sb_2__2__13_chanx_right_out;
wire [0:95] sb_2__2__13_chany_bottom_out;
wire [0:95] sb_2__2__13_chany_top_out;
wire [0:95] sb_2__2__14_chanx_left_out;
wire [0:95] sb_2__2__14_chanx_right_out;
wire [0:95] sb_2__2__14_chany_bottom_out;
wire [0:95] sb_2__2__14_chany_top_out;
wire [0:95] sb_2__2__1_chanx_left_out;
wire [0:95] sb_2__2__1_chanx_right_out;
wire [0:95] sb_2__2__1_chany_bottom_out;
wire [0:95] sb_2__2__1_chany_top_out;
wire [0:95] sb_2__2__2_chanx_left_out;
wire [0:95] sb_2__2__2_chanx_right_out;
wire [0:95] sb_2__2__2_chany_bottom_out;
wire [0:95] sb_2__2__2_chany_top_out;
wire [0:95] sb_2__2__3_chanx_left_out;
wire [0:95] sb_2__2__3_chanx_right_out;
wire [0:95] sb_2__2__3_chany_bottom_out;
wire [0:95] sb_2__2__3_chany_top_out;
wire [0:95] sb_2__2__4_chanx_left_out;
wire [0:95] sb_2__2__4_chanx_right_out;
wire [0:95] sb_2__2__4_chany_bottom_out;
wire [0:95] sb_2__2__4_chany_top_out;
wire [0:95] sb_2__2__5_chanx_left_out;
wire [0:95] sb_2__2__5_chanx_right_out;
wire [0:95] sb_2__2__5_chany_bottom_out;
wire [0:95] sb_2__2__5_chany_top_out;
wire [0:95] sb_2__2__6_chanx_left_out;
wire [0:95] sb_2__2__6_chanx_right_out;
wire [0:95] sb_2__2__6_chany_bottom_out;
wire [0:95] sb_2__2__6_chany_top_out;
wire [0:95] sb_2__2__7_chanx_left_out;
wire [0:95] sb_2__2__7_chanx_right_out;
wire [0:95] sb_2__2__7_chany_bottom_out;
wire [0:95] sb_2__2__7_chany_top_out;
wire [0:95] sb_2__2__8_chanx_left_out;
wire [0:95] sb_2__2__8_chanx_right_out;
wire [0:95] sb_2__2__8_chany_bottom_out;
wire [0:95] sb_2__2__8_chany_top_out;
wire [0:95] sb_2__2__9_chanx_left_out;
wire [0:95] sb_2__2__9_chanx_right_out;
wire [0:95] sb_2__2__9_chany_bottom_out;
wire [0:95] sb_2__2__9_chany_top_out;
wire [0:95] sb_2__7__0_chanx_left_out;
wire [0:95] sb_2__7__0_chanx_right_out;
wire [0:95] sb_2__7__0_chany_bottom_out;
wire [0:95] sb_2__7__0_chany_top_out;
wire [0:95] sb_2__7__1_chanx_left_out;
wire [0:95] sb_2__7__1_chanx_right_out;
wire [0:95] sb_2__7__1_chany_bottom_out;
wire [0:95] sb_2__7__1_chany_top_out;
wire [0:95] sb_2__7__2_chanx_left_out;
wire [0:95] sb_2__7__2_chanx_right_out;
wire [0:95] sb_2__7__2_chany_bottom_out;
wire [0:95] sb_2__7__2_chany_top_out;
wire [0:95] sb_2__8__0_chanx_left_out;
wire [0:95] sb_2__8__0_chanx_right_out;
wire [0:95] sb_2__8__0_chany_bottom_out;
wire [0:95] sb_2__8__1_chanx_left_out;
wire [0:95] sb_2__8__1_chanx_right_out;
wire [0:95] sb_2__8__1_chany_bottom_out;
wire [0:95] sb_2__8__2_chanx_left_out;
wire [0:95] sb_2__8__2_chanx_right_out;
wire [0:95] sb_2__8__2_chany_bottom_out;
wire [0:95] sb_2__8__3_chanx_left_out;
wire [0:95] sb_2__8__3_chanx_right_out;
wire [0:95] sb_2__8__3_chany_bottom_out;
wire [0:95] sb_2__8__4_chanx_left_out;
wire [0:95] sb_2__8__4_chanx_right_out;
wire [0:95] sb_2__8__4_chany_bottom_out;
wire [0:95] sb_2__8__5_chanx_left_out;
wire [0:95] sb_2__8__5_chanx_right_out;
wire [0:95] sb_2__8__5_chany_bottom_out;
wire [0:95] sb_2__8__6_chanx_left_out;
wire [0:95] sb_2__8__6_chanx_right_out;
wire [0:95] sb_2__8__6_chany_bottom_out;
wire [0:95] sb_3__1__0_chanx_left_out;
wire [0:95] sb_3__1__0_chanx_right_out;
wire [0:95] sb_3__1__0_chany_bottom_out;
wire [0:95] sb_3__1__0_chany_top_out;
wire [0:95] sb_3__2__0_chanx_left_out;
wire [0:95] sb_3__2__0_chanx_right_out;
wire [0:95] sb_3__2__0_chany_bottom_out;
wire [0:95] sb_3__2__0_chany_top_out;
wire [0:95] sb_3__2__1_chanx_left_out;
wire [0:95] sb_3__2__1_chanx_right_out;
wire [0:95] sb_3__2__1_chany_bottom_out;
wire [0:95] sb_3__2__1_chany_top_out;
wire [0:95] sb_3__2__2_chanx_left_out;
wire [0:95] sb_3__2__2_chanx_right_out;
wire [0:95] sb_3__2__2_chany_bottom_out;
wire [0:95] sb_3__2__2_chany_top_out;
wire [0:95] sb_3__2__3_chanx_left_out;
wire [0:95] sb_3__2__3_chanx_right_out;
wire [0:95] sb_3__2__3_chany_bottom_out;
wire [0:95] sb_3__2__3_chany_top_out;
wire [0:95] sb_3__2__4_chanx_left_out;
wire [0:95] sb_3__2__4_chanx_right_out;
wire [0:95] sb_3__2__4_chany_bottom_out;
wire [0:95] sb_3__2__4_chany_top_out;
wire [0:95] sb_3__2__5_chanx_left_out;
wire [0:95] sb_3__2__5_chanx_right_out;
wire [0:95] sb_3__2__5_chany_bottom_out;
wire [0:95] sb_3__2__5_chany_top_out;
wire [0:95] sb_3__2__6_chanx_left_out;
wire [0:95] sb_3__2__6_chanx_right_out;
wire [0:95] sb_3__2__6_chany_bottom_out;
wire [0:95] sb_3__2__6_chany_top_out;
wire [0:95] sb_3__2__7_chanx_left_out;
wire [0:95] sb_3__2__7_chanx_right_out;
wire [0:95] sb_3__2__7_chany_bottom_out;
wire [0:95] sb_3__2__7_chany_top_out;
wire [0:95] sb_3__2__8_chanx_left_out;
wire [0:95] sb_3__2__8_chanx_right_out;
wire [0:95] sb_3__2__8_chany_bottom_out;
wire [0:95] sb_3__2__8_chany_top_out;
wire [0:95] sb_3__4__0_chanx_left_out;
wire [0:95] sb_3__4__0_chanx_right_out;
wire [0:95] sb_3__4__0_chany_bottom_out;
wire [0:95] sb_3__4__0_chany_top_out;
wire [0:95] sb_3__7__0_chanx_left_out;
wire [0:95] sb_3__7__0_chanx_right_out;
wire [0:95] sb_3__7__0_chany_bottom_out;
wire [0:95] sb_3__7__0_chany_top_out;
wire [0:95] sb_3__7__1_chanx_left_out;
wire [0:95] sb_3__7__1_chanx_right_out;
wire [0:95] sb_3__7__1_chany_bottom_out;
wire [0:95] sb_3__7__1_chany_top_out;
wire [0:95] sb_4__1__0_chanx_left_out;
wire [0:95] sb_4__1__0_chanx_right_out;
wire [0:95] sb_4__1__0_chany_bottom_out;
wire [0:95] sb_4__1__0_chany_top_out;
wire [0:95] sb_4__2__0_chanx_left_out;
wire [0:95] sb_4__2__0_chanx_right_out;
wire [0:95] sb_4__2__0_chany_bottom_out;
wire [0:95] sb_4__2__0_chany_top_out;
wire [0:95] sb_4__2__1_chanx_left_out;
wire [0:95] sb_4__2__1_chanx_right_out;
wire [0:95] sb_4__2__1_chany_bottom_out;
wire [0:95] sb_4__2__1_chany_top_out;
wire [0:95] sb_4__3__0_chanx_left_out;
wire [0:95] sb_4__3__0_chanx_right_out;
wire [0:95] sb_4__3__0_chany_bottom_out;
wire [0:95] sb_4__3__0_chany_top_out;
wire [0:95] sb_4__3__1_chanx_left_out;
wire [0:95] sb_4__3__1_chanx_right_out;
wire [0:95] sb_4__3__1_chany_bottom_out;
wire [0:95] sb_4__3__1_chany_top_out;
wire [0:95] sb_4__4__0_chanx_left_out;
wire [0:95] sb_4__4__0_chanx_right_out;
wire [0:95] sb_4__4__0_chany_bottom_out;
wire [0:95] sb_4__4__0_chany_top_out;
wire [0:95] sb_4__7__0_chanx_left_out;
wire [0:95] sb_4__7__0_chanx_right_out;
wire [0:95] sb_4__7__0_chany_bottom_out;
wire [0:95] sb_4__7__0_chany_top_out;
wire [0:95] sb_7__1__0_chanx_left_out;
wire [0:95] sb_7__1__0_chanx_right_out;
wire [0:95] sb_7__1__0_chany_bottom_out;
wire [0:95] sb_7__1__0_chany_top_out;
wire [0:95] sb_7__2__0_chanx_left_out;
wire [0:95] sb_7__2__0_chanx_right_out;
wire [0:95] sb_7__2__0_chany_bottom_out;
wire [0:95] sb_7__2__0_chany_top_out;
wire [0:95] sb_7__2__1_chanx_left_out;
wire [0:95] sb_7__2__1_chanx_right_out;
wire [0:95] sb_7__2__1_chany_bottom_out;
wire [0:95] sb_7__2__1_chany_top_out;
wire [0:95] sb_7__2__2_chanx_left_out;
wire [0:95] sb_7__2__2_chanx_right_out;
wire [0:95] sb_7__2__2_chany_bottom_out;
wire [0:95] sb_7__2__2_chany_top_out;
wire [0:95] sb_7__2__3_chanx_left_out;
wire [0:95] sb_7__2__3_chanx_right_out;
wire [0:95] sb_7__2__3_chany_bottom_out;
wire [0:95] sb_7__2__3_chany_top_out;
wire [0:95] sb_7__2__4_chanx_left_out;
wire [0:95] sb_7__2__4_chanx_right_out;
wire [0:95] sb_7__2__4_chany_bottom_out;
wire [0:95] sb_7__2__4_chany_top_out;
wire [0:95] sb_7__7__0_chanx_left_out;
wire [0:95] sb_7__7__0_chanx_right_out;
wire [0:95] sb_7__7__0_chany_bottom_out;
wire [0:95] sb_7__7__0_chany_top_out;
wire [0:95] sb_9__1__0_chanx_left_out;
wire [0:95] sb_9__1__0_chanx_right_out;
wire [0:95] sb_9__1__0_chany_bottom_out;
wire [0:95] sb_9__1__0_chany_top_out;
wire [0:95] sb_9__2__0_chanx_left_out;
wire [0:95] sb_9__2__0_chanx_right_out;
wire [0:95] sb_9__2__0_chany_bottom_out;
wire [0:95] sb_9__2__0_chany_top_out;
wire [0:95] sb_9__2__1_chanx_left_out;
wire [0:95] sb_9__2__1_chanx_right_out;
wire [0:95] sb_9__2__1_chany_bottom_out;
wire [0:95] sb_9__2__1_chany_top_out;
wire [0:95] sb_9__2__2_chanx_left_out;
wire [0:95] sb_9__2__2_chanx_right_out;
wire [0:95] sb_9__2__2_chany_bottom_out;
wire [0:95] sb_9__2__2_chany_top_out;
wire [0:95] sb_9__2__3_chanx_left_out;
wire [0:95] sb_9__2__3_chanx_right_out;
wire [0:95] sb_9__2__3_chany_bottom_out;
wire [0:95] sb_9__2__3_chany_top_out;
wire [0:95] sb_9__2__4_chanx_left_out;
wire [0:95] sb_9__2__4_chanx_right_out;
wire [0:95] sb_9__2__4_chany_bottom_out;
wire [0:95] sb_9__2__4_chany_top_out;
wire [0:95] sb_9__7__0_chanx_left_out;
wire [0:95] sb_9__7__0_chanx_right_out;
wire [0:95] sb_9__7__0_chany_bottom_out;
wire [0:95] sb_9__7__0_chany_top_out;

// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	grid_io_left grid_io_left_1__1_ (
		.test_en(test_en),
		.scan_mode(scan_mode),
		.scan_clk(scan_clk),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.CFG_DONE(CFG_DONE),
		.gfpga_pad_QL_PREIO_A2F(gfpga_pad_QL_PREIO_A2F[0:19]),
		.gfpga_pad_QL_PREIO_F2A(gfpga_pad_QL_PREIO_F2A[0:19]),
		.gfpga_pad_QL_PREIO_F2A_DEF0(gfpga_pad_QL_PREIO_F2A_DEF0[0:19]),
		.gfpga_pad_QL_PREIO_F2A_DEF1(gfpga_pad_QL_PREIO_F2A_DEF1[0:19]),
		.gfpga_pad_QL_PREIO_F2A_CLK(gfpga_pad_QL_PREIO_F2A_CLK[0:19]),
		.right_width_0_height_0_subtile_0__pin_f2a_i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_0__pin_sc_in_0_(grid_io_left_1__1__undriven_right_width_0_height_0_subtile_0__pin_sc_in_0_),
		.right_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_1__pin_f2a_i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_1__pin_sc_in_0_(grid_io_left_1__1__undriven_right_width_0_height_0_subtile_1__pin_sc_in_0_),
		.right_width_0_height_0_subtile_1__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_1__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_1__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_1__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_1__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_1__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_2__pin_f2a_i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_2__pin_sc_in_0_(grid_io_left_1__1__undriven_right_width_0_height_0_subtile_2__pin_sc_in_0_),
		.right_width_0_height_0_subtile_2__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_2__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_2__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_2__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_2__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_2__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_3__pin_f2a_i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_3__pin_sc_in_0_(grid_io_left_1__1__undriven_right_width_0_height_0_subtile_3__pin_sc_in_0_),
		.right_width_0_height_0_subtile_3__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_3__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_3__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_3__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_3__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_3__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_4__pin_f2a_i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_4__pin_sc_in_0_(grid_io_left_1__1__undriven_right_width_0_height_0_subtile_4__pin_sc_in_0_),
		.right_width_0_height_0_subtile_4__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_4__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_4__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_4__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_4__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_4__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_5__pin_f2a_i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_5__pin_sc_in_0_(grid_io_left_1__1__undriven_right_width_0_height_0_subtile_5__pin_sc_in_0_),
		.right_width_0_height_0_subtile_5__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_5__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_5__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_5__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_5__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_5__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_6__pin_f2a_i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_6__pin_sc_in_0_(grid_io_left_1__1__undriven_right_width_0_height_0_subtile_6__pin_sc_in_0_),
		.right_width_0_height_0_subtile_6__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_6__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_6__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_6__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_6__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_6__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_7__pin_f2a_i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_7__pin_sc_in_0_(grid_io_left_1__1__undriven_right_width_0_height_0_subtile_7__pin_sc_in_0_),
		.right_width_0_height_0_subtile_7__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_7__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_7__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_7__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_7__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_7__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_8__pin_f2a_i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_8__pin_sc_in_0_(grid_io_left_1__1__undriven_right_width_0_height_0_subtile_8__pin_sc_in_0_),
		.right_width_0_height_0_subtile_8__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_8__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_8__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_8__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_8__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_8__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_9__pin_f2a_i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_9__pin_sc_in_0_(grid_io_left_1__1__undriven_right_width_0_height_0_subtile_9__pin_sc_in_0_),
		.right_width_0_height_0_subtile_9__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_9__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_9__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_9__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_9__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_9__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_10__pin_f2a_i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_10__pin_sc_in_0_(grid_io_left_1__1__undriven_right_width_0_height_0_subtile_10__pin_sc_in_0_),
		.right_width_0_height_0_subtile_10__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_10__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_10__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_10__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_10__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_10__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_11__pin_f2a_i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_11__pin_sc_in_0_(grid_io_left_1__1__undriven_right_width_0_height_0_subtile_11__pin_sc_in_0_),
		.right_width_0_height_0_subtile_11__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_11__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_11__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_11__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_11__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_11__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_12__pin_f2a_i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_12__pin_sc_in_0_(grid_io_left_1__1__undriven_right_width_0_height_0_subtile_12__pin_sc_in_0_),
		.right_width_0_height_0_subtile_12__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_12__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_12__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_12__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_12__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_12__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_13__pin_f2a_i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_13__pin_sc_in_0_(grid_io_left_1__1__undriven_right_width_0_height_0_subtile_13__pin_sc_in_0_),
		.right_width_0_height_0_subtile_13__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_13__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_13__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_13__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_13__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_13__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_14__pin_f2a_i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_14__pin_sc_in_0_(grid_io_left_1__1__undriven_right_width_0_height_0_subtile_14__pin_sc_in_0_),
		.right_width_0_height_0_subtile_14__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_14__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_14__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_14__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_14__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_14__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_15__pin_f2a_i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_15__pin_sc_in_0_(grid_io_left_1__1__undriven_right_width_0_height_0_subtile_15__pin_sc_in_0_),
		.right_width_0_height_0_subtile_15__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_15__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_15__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_15__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_15__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_15__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_16__pin_f2a_i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_16__pin_sc_in_0_(grid_io_left_1__1__undriven_right_width_0_height_0_subtile_16__pin_sc_in_0_),
		.right_width_0_height_0_subtile_16__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_16__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_16__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_16__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_16__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_16__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_17__pin_f2a_i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_17__pin_sc_in_0_(grid_io_left_1__1__undriven_right_width_0_height_0_subtile_17__pin_sc_in_0_),
		.right_width_0_height_0_subtile_17__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_17__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_17__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_17__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_17__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_17__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_18__pin_f2a_i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_18__pin_sc_in_0_(grid_io_left_1__1__undriven_right_width_0_height_0_subtile_18__pin_sc_in_0_),
		.right_width_0_height_0_subtile_18__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_18__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_18__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_18__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_18__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_18__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_19__pin_f2a_i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_19__pin_sc_in_0_(grid_io_left_1__1__undriven_right_width_0_height_0_subtile_19__pin_sc_in_0_),
		.right_width_0_height_0_subtile_19__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_19__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_19__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_19__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_19__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_19__pin_clk_3_(clk[3]),
		.ccff_head(cby_1__1__0_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_0__pin_sc_out_0_(grid_io_left_1__1__undriven_right_width_0_height_0_subtile_0__pin_sc_out_0_),
		.right_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_1__pin_sc_out_0_(grid_io_left_1__1__undriven_right_width_0_height_0_subtile_1__pin_sc_out_0_),
		.right_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_2__pin_sc_out_0_(grid_io_left_1__1__undriven_right_width_0_height_0_subtile_2__pin_sc_out_0_),
		.right_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_3__pin_sc_out_0_(grid_io_left_1__1__undriven_right_width_0_height_0_subtile_3__pin_sc_out_0_),
		.right_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_4__pin_sc_out_0_(grid_io_left_1__1__undriven_right_width_0_height_0_subtile_4__pin_sc_out_0_),
		.right_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_5__pin_sc_out_0_(grid_io_left_1__1__undriven_right_width_0_height_0_subtile_5__pin_sc_out_0_),
		.right_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_6__pin_sc_out_0_(grid_io_left_1__1__undriven_right_width_0_height_0_subtile_6__pin_sc_out_0_),
		.right_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_7__pin_sc_out_0_(grid_io_left_1__1__undriven_right_width_0_height_0_subtile_7__pin_sc_out_0_),
		.right_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_8__pin_sc_out_0_(grid_io_left_1__1__undriven_right_width_0_height_0_subtile_8__pin_sc_out_0_),
		.right_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_9__pin_sc_out_0_(grid_io_left_1__1__undriven_right_width_0_height_0_subtile_9__pin_sc_out_0_),
		.right_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_10__pin_sc_out_0_(grid_io_left_1__1__undriven_right_width_0_height_0_subtile_10__pin_sc_out_0_),
		.right_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_11__pin_sc_out_0_(grid_io_left_1__1__undriven_right_width_0_height_0_subtile_11__pin_sc_out_0_),
		.right_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_12__pin_sc_out_0_(grid_io_left_1__1__undriven_right_width_0_height_0_subtile_12__pin_sc_out_0_),
		.right_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_13__pin_sc_out_0_(grid_io_left_1__1__undriven_right_width_0_height_0_subtile_13__pin_sc_out_0_),
		.right_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_14__pin_sc_out_0_(grid_io_left_1__1__undriven_right_width_0_height_0_subtile_14__pin_sc_out_0_),
		.right_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_15__pin_sc_out_0_(grid_io_left_1__1__undriven_right_width_0_height_0_subtile_15__pin_sc_out_0_),
		.right_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_16__pin_sc_out_0_(grid_io_left_1__1__undriven_right_width_0_height_0_subtile_16__pin_sc_out_0_),
		.right_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_17__pin_sc_out_0_(grid_io_left_1__1__undriven_right_width_0_height_0_subtile_17__pin_sc_out_0_),
		.right_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_18__pin_sc_out_0_(grid_io_left_1__1__undriven_right_width_0_height_0_subtile_18__pin_sc_out_0_),
		.right_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_19__pin_sc_out_0_(grid_io_left_1__1__undriven_right_width_0_height_0_subtile_19__pin_sc_out_0_),
		.ccff_tail(grid_io_left_0_ccff_tail));

	grid_io_left grid_io_left_1__2_ (
		.test_en(test_en),
		.scan_mode(scan_mode),
		.scan_clk(scan_clk),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.CFG_DONE(CFG_DONE),
		.gfpga_pad_QL_PREIO_A2F(gfpga_pad_QL_PREIO_A2F[20:39]),
		.gfpga_pad_QL_PREIO_F2A(gfpga_pad_QL_PREIO_F2A[20:39]),
		.gfpga_pad_QL_PREIO_F2A_DEF0(gfpga_pad_QL_PREIO_F2A_DEF0[20:39]),
		.gfpga_pad_QL_PREIO_F2A_DEF1(gfpga_pad_QL_PREIO_F2A_DEF1[20:39]),
		.gfpga_pad_QL_PREIO_F2A_CLK(gfpga_pad_QL_PREIO_F2A_CLK[20:39]),
		.right_width_0_height_0_subtile_0__pin_f2a_i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_0__pin_sc_in_0_(grid_io_left_1__2__undriven_right_width_0_height_0_subtile_0__pin_sc_in_0_),
		.right_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_1__pin_f2a_i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_1__pin_sc_in_0_(grid_io_left_1__2__undriven_right_width_0_height_0_subtile_1__pin_sc_in_0_),
		.right_width_0_height_0_subtile_1__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_1__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_1__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_1__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_1__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_1__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_2__pin_f2a_i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_2__pin_sc_in_0_(grid_io_left_1__2__undriven_right_width_0_height_0_subtile_2__pin_sc_in_0_),
		.right_width_0_height_0_subtile_2__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_2__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_2__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_2__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_2__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_2__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_3__pin_f2a_i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_3__pin_sc_in_0_(grid_io_left_1__2__undriven_right_width_0_height_0_subtile_3__pin_sc_in_0_),
		.right_width_0_height_0_subtile_3__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_3__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_3__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_3__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_3__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_3__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_4__pin_f2a_i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_4__pin_sc_in_0_(grid_io_left_1__2__undriven_right_width_0_height_0_subtile_4__pin_sc_in_0_),
		.right_width_0_height_0_subtile_4__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_4__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_4__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_4__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_4__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_4__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_5__pin_f2a_i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_5__pin_sc_in_0_(grid_io_left_1__2__undriven_right_width_0_height_0_subtile_5__pin_sc_in_0_),
		.right_width_0_height_0_subtile_5__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_5__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_5__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_5__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_5__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_5__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_6__pin_f2a_i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_6__pin_sc_in_0_(grid_io_left_1__2__undriven_right_width_0_height_0_subtile_6__pin_sc_in_0_),
		.right_width_0_height_0_subtile_6__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_6__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_6__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_6__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_6__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_6__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_7__pin_f2a_i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_7__pin_sc_in_0_(grid_io_left_1__2__undriven_right_width_0_height_0_subtile_7__pin_sc_in_0_),
		.right_width_0_height_0_subtile_7__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_7__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_7__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_7__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_7__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_7__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_8__pin_f2a_i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_8__pin_sc_in_0_(grid_io_left_1__2__undriven_right_width_0_height_0_subtile_8__pin_sc_in_0_),
		.right_width_0_height_0_subtile_8__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_8__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_8__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_8__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_8__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_8__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_9__pin_f2a_i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_9__pin_sc_in_0_(grid_io_left_1__2__undriven_right_width_0_height_0_subtile_9__pin_sc_in_0_),
		.right_width_0_height_0_subtile_9__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_9__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_9__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_9__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_9__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_9__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_10__pin_f2a_i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_10__pin_sc_in_0_(grid_io_left_1__2__undriven_right_width_0_height_0_subtile_10__pin_sc_in_0_),
		.right_width_0_height_0_subtile_10__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_10__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_10__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_10__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_10__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_10__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_11__pin_f2a_i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_11__pin_sc_in_0_(grid_io_left_1__2__undriven_right_width_0_height_0_subtile_11__pin_sc_in_0_),
		.right_width_0_height_0_subtile_11__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_11__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_11__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_11__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_11__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_11__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_12__pin_f2a_i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_12__pin_sc_in_0_(grid_io_left_1__2__undriven_right_width_0_height_0_subtile_12__pin_sc_in_0_),
		.right_width_0_height_0_subtile_12__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_12__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_12__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_12__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_12__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_12__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_13__pin_f2a_i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_13__pin_sc_in_0_(grid_io_left_1__2__undriven_right_width_0_height_0_subtile_13__pin_sc_in_0_),
		.right_width_0_height_0_subtile_13__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_13__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_13__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_13__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_13__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_13__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_14__pin_f2a_i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_14__pin_sc_in_0_(grid_io_left_1__2__undriven_right_width_0_height_0_subtile_14__pin_sc_in_0_),
		.right_width_0_height_0_subtile_14__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_14__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_14__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_14__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_14__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_14__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_15__pin_f2a_i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_15__pin_sc_in_0_(grid_io_left_1__2__undriven_right_width_0_height_0_subtile_15__pin_sc_in_0_),
		.right_width_0_height_0_subtile_15__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_15__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_15__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_15__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_15__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_15__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_16__pin_f2a_i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_16__pin_sc_in_0_(grid_io_left_1__2__undriven_right_width_0_height_0_subtile_16__pin_sc_in_0_),
		.right_width_0_height_0_subtile_16__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_16__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_16__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_16__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_16__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_16__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_17__pin_f2a_i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_17__pin_sc_in_0_(grid_io_left_1__2__undriven_right_width_0_height_0_subtile_17__pin_sc_in_0_),
		.right_width_0_height_0_subtile_17__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_17__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_17__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_17__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_17__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_17__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_18__pin_f2a_i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_18__pin_sc_in_0_(grid_io_left_1__2__undriven_right_width_0_height_0_subtile_18__pin_sc_in_0_),
		.right_width_0_height_0_subtile_18__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_18__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_18__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_18__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_18__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_18__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_19__pin_f2a_i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_19__pin_sc_in_0_(grid_io_left_1__2__undriven_right_width_0_height_0_subtile_19__pin_sc_in_0_),
		.right_width_0_height_0_subtile_19__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_19__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_19__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_19__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_19__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_19__pin_clk_3_(clk[3]),
		.ccff_head(cby_1__1__1_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_0__pin_sc_out_0_(grid_io_left_1__2__undriven_right_width_0_height_0_subtile_0__pin_sc_out_0_),
		.right_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_1__pin_sc_out_0_(grid_io_left_1__2__undriven_right_width_0_height_0_subtile_1__pin_sc_out_0_),
		.right_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_2__pin_sc_out_0_(grid_io_left_1__2__undriven_right_width_0_height_0_subtile_2__pin_sc_out_0_),
		.right_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_3__pin_sc_out_0_(grid_io_left_1__2__undriven_right_width_0_height_0_subtile_3__pin_sc_out_0_),
		.right_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_4__pin_sc_out_0_(grid_io_left_1__2__undriven_right_width_0_height_0_subtile_4__pin_sc_out_0_),
		.right_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_5__pin_sc_out_0_(grid_io_left_1__2__undriven_right_width_0_height_0_subtile_5__pin_sc_out_0_),
		.right_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_6__pin_sc_out_0_(grid_io_left_1__2__undriven_right_width_0_height_0_subtile_6__pin_sc_out_0_),
		.right_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_7__pin_sc_out_0_(grid_io_left_1__2__undriven_right_width_0_height_0_subtile_7__pin_sc_out_0_),
		.right_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_8__pin_sc_out_0_(grid_io_left_1__2__undriven_right_width_0_height_0_subtile_8__pin_sc_out_0_),
		.right_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_9__pin_sc_out_0_(grid_io_left_1__2__undriven_right_width_0_height_0_subtile_9__pin_sc_out_0_),
		.right_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_10__pin_sc_out_0_(grid_io_left_1__2__undriven_right_width_0_height_0_subtile_10__pin_sc_out_0_),
		.right_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_11__pin_sc_out_0_(grid_io_left_1__2__undriven_right_width_0_height_0_subtile_11__pin_sc_out_0_),
		.right_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_12__pin_sc_out_0_(grid_io_left_1__2__undriven_right_width_0_height_0_subtile_12__pin_sc_out_0_),
		.right_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_13__pin_sc_out_0_(grid_io_left_1__2__undriven_right_width_0_height_0_subtile_13__pin_sc_out_0_),
		.right_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_14__pin_sc_out_0_(grid_io_left_1__2__undriven_right_width_0_height_0_subtile_14__pin_sc_out_0_),
		.right_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_15__pin_sc_out_0_(grid_io_left_1__2__undriven_right_width_0_height_0_subtile_15__pin_sc_out_0_),
		.right_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_16__pin_sc_out_0_(grid_io_left_1__2__undriven_right_width_0_height_0_subtile_16__pin_sc_out_0_),
		.right_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_17__pin_sc_out_0_(grid_io_left_1__2__undriven_right_width_0_height_0_subtile_17__pin_sc_out_0_),
		.right_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_18__pin_sc_out_0_(grid_io_left_1__2__undriven_right_width_0_height_0_subtile_18__pin_sc_out_0_),
		.right_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_19__pin_sc_out_0_(grid_io_left_1__2__undriven_right_width_0_height_0_subtile_19__pin_sc_out_0_),
		.ccff_tail(grid_io_left_1_ccff_tail));

	grid_io_left grid_io_left_1__3_ (
		.test_en(test_en),
		.scan_mode(scan_mode),
		.scan_clk(scan_clk),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.CFG_DONE(CFG_DONE),
		.gfpga_pad_QL_PREIO_A2F(gfpga_pad_QL_PREIO_A2F[40:59]),
		.gfpga_pad_QL_PREIO_F2A(gfpga_pad_QL_PREIO_F2A[40:59]),
		.gfpga_pad_QL_PREIO_F2A_DEF0(gfpga_pad_QL_PREIO_F2A_DEF0[40:59]),
		.gfpga_pad_QL_PREIO_F2A_DEF1(gfpga_pad_QL_PREIO_F2A_DEF1[40:59]),
		.gfpga_pad_QL_PREIO_F2A_CLK(gfpga_pad_QL_PREIO_F2A_CLK[40:59]),
		.right_width_0_height_0_subtile_0__pin_f2a_i_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_0__pin_sc_in_0_(grid_io_left_1__3__undriven_right_width_0_height_0_subtile_0__pin_sc_in_0_),
		.right_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_1__pin_f2a_i_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_1__pin_sc_in_0_(grid_io_left_1__3__undriven_right_width_0_height_0_subtile_1__pin_sc_in_0_),
		.right_width_0_height_0_subtile_1__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_1__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_1__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_1__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_1__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_1__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_2__pin_f2a_i_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_2__pin_sc_in_0_(grid_io_left_1__3__undriven_right_width_0_height_0_subtile_2__pin_sc_in_0_),
		.right_width_0_height_0_subtile_2__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_2__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_2__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_2__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_2__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_2__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_3__pin_f2a_i_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_3__pin_sc_in_0_(grid_io_left_1__3__undriven_right_width_0_height_0_subtile_3__pin_sc_in_0_),
		.right_width_0_height_0_subtile_3__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_3__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_3__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_3__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_3__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_3__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_4__pin_f2a_i_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_4__pin_sc_in_0_(grid_io_left_1__3__undriven_right_width_0_height_0_subtile_4__pin_sc_in_0_),
		.right_width_0_height_0_subtile_4__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_4__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_4__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_4__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_4__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_4__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_5__pin_f2a_i_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_5__pin_sc_in_0_(grid_io_left_1__3__undriven_right_width_0_height_0_subtile_5__pin_sc_in_0_),
		.right_width_0_height_0_subtile_5__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_5__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_5__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_5__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_5__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_5__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_6__pin_f2a_i_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_6__pin_sc_in_0_(grid_io_left_1__3__undriven_right_width_0_height_0_subtile_6__pin_sc_in_0_),
		.right_width_0_height_0_subtile_6__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_6__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_6__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_6__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_6__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_6__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_7__pin_f2a_i_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_7__pin_sc_in_0_(grid_io_left_1__3__undriven_right_width_0_height_0_subtile_7__pin_sc_in_0_),
		.right_width_0_height_0_subtile_7__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_7__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_7__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_7__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_7__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_7__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_8__pin_f2a_i_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_8__pin_sc_in_0_(grid_io_left_1__3__undriven_right_width_0_height_0_subtile_8__pin_sc_in_0_),
		.right_width_0_height_0_subtile_8__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_8__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_8__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_8__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_8__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_8__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_9__pin_f2a_i_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_9__pin_sc_in_0_(grid_io_left_1__3__undriven_right_width_0_height_0_subtile_9__pin_sc_in_0_),
		.right_width_0_height_0_subtile_9__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_9__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_9__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_9__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_9__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_9__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_10__pin_f2a_i_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_10__pin_sc_in_0_(grid_io_left_1__3__undriven_right_width_0_height_0_subtile_10__pin_sc_in_0_),
		.right_width_0_height_0_subtile_10__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_10__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_10__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_10__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_10__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_10__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_11__pin_f2a_i_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_11__pin_sc_in_0_(grid_io_left_1__3__undriven_right_width_0_height_0_subtile_11__pin_sc_in_0_),
		.right_width_0_height_0_subtile_11__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_11__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_11__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_11__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_11__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_11__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_12__pin_f2a_i_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_12__pin_sc_in_0_(grid_io_left_1__3__undriven_right_width_0_height_0_subtile_12__pin_sc_in_0_),
		.right_width_0_height_0_subtile_12__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_12__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_12__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_12__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_12__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_12__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_13__pin_f2a_i_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_13__pin_sc_in_0_(grid_io_left_1__3__undriven_right_width_0_height_0_subtile_13__pin_sc_in_0_),
		.right_width_0_height_0_subtile_13__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_13__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_13__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_13__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_13__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_13__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_14__pin_f2a_i_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_14__pin_sc_in_0_(grid_io_left_1__3__undriven_right_width_0_height_0_subtile_14__pin_sc_in_0_),
		.right_width_0_height_0_subtile_14__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_14__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_14__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_14__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_14__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_14__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_15__pin_f2a_i_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_15__pin_sc_in_0_(grid_io_left_1__3__undriven_right_width_0_height_0_subtile_15__pin_sc_in_0_),
		.right_width_0_height_0_subtile_15__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_15__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_15__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_15__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_15__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_15__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_16__pin_f2a_i_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_16__pin_sc_in_0_(grid_io_left_1__3__undriven_right_width_0_height_0_subtile_16__pin_sc_in_0_),
		.right_width_0_height_0_subtile_16__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_16__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_16__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_16__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_16__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_16__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_17__pin_f2a_i_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_17__pin_sc_in_0_(grid_io_left_1__3__undriven_right_width_0_height_0_subtile_17__pin_sc_in_0_),
		.right_width_0_height_0_subtile_17__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_17__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_17__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_17__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_17__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_17__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_18__pin_f2a_i_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_18__pin_sc_in_0_(grid_io_left_1__3__undriven_right_width_0_height_0_subtile_18__pin_sc_in_0_),
		.right_width_0_height_0_subtile_18__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_18__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_18__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_18__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_18__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_18__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_19__pin_f2a_i_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_19__pin_sc_in_0_(grid_io_left_1__3__undriven_right_width_0_height_0_subtile_19__pin_sc_in_0_),
		.right_width_0_height_0_subtile_19__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_19__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_19__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_19__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_19__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_19__pin_clk_3_(clk[3]),
		.ccff_head(cby_1__1__2_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_0__pin_sc_out_0_(grid_io_left_1__3__undriven_right_width_0_height_0_subtile_0__pin_sc_out_0_),
		.right_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_1__pin_sc_out_0_(grid_io_left_1__3__undriven_right_width_0_height_0_subtile_1__pin_sc_out_0_),
		.right_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_2__pin_sc_out_0_(grid_io_left_1__3__undriven_right_width_0_height_0_subtile_2__pin_sc_out_0_),
		.right_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_3__pin_sc_out_0_(grid_io_left_1__3__undriven_right_width_0_height_0_subtile_3__pin_sc_out_0_),
		.right_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_4__pin_sc_out_0_(grid_io_left_1__3__undriven_right_width_0_height_0_subtile_4__pin_sc_out_0_),
		.right_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_5__pin_sc_out_0_(grid_io_left_1__3__undriven_right_width_0_height_0_subtile_5__pin_sc_out_0_),
		.right_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_6__pin_sc_out_0_(grid_io_left_1__3__undriven_right_width_0_height_0_subtile_6__pin_sc_out_0_),
		.right_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_7__pin_sc_out_0_(grid_io_left_1__3__undriven_right_width_0_height_0_subtile_7__pin_sc_out_0_),
		.right_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_8__pin_sc_out_0_(grid_io_left_1__3__undriven_right_width_0_height_0_subtile_8__pin_sc_out_0_),
		.right_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_9__pin_sc_out_0_(grid_io_left_1__3__undriven_right_width_0_height_0_subtile_9__pin_sc_out_0_),
		.right_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_10__pin_sc_out_0_(grid_io_left_1__3__undriven_right_width_0_height_0_subtile_10__pin_sc_out_0_),
		.right_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_11__pin_sc_out_0_(grid_io_left_1__3__undriven_right_width_0_height_0_subtile_11__pin_sc_out_0_),
		.right_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_12__pin_sc_out_0_(grid_io_left_1__3__undriven_right_width_0_height_0_subtile_12__pin_sc_out_0_),
		.right_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_13__pin_sc_out_0_(grid_io_left_1__3__undriven_right_width_0_height_0_subtile_13__pin_sc_out_0_),
		.right_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_14__pin_sc_out_0_(grid_io_left_1__3__undriven_right_width_0_height_0_subtile_14__pin_sc_out_0_),
		.right_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_15__pin_sc_out_0_(grid_io_left_1__3__undriven_right_width_0_height_0_subtile_15__pin_sc_out_0_),
		.right_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_16__pin_sc_out_0_(grid_io_left_1__3__undriven_right_width_0_height_0_subtile_16__pin_sc_out_0_),
		.right_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_17__pin_sc_out_0_(grid_io_left_1__3__undriven_right_width_0_height_0_subtile_17__pin_sc_out_0_),
		.right_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_18__pin_sc_out_0_(grid_io_left_1__3__undriven_right_width_0_height_0_subtile_18__pin_sc_out_0_),
		.right_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_19__pin_sc_out_0_(grid_io_left_1__3__undriven_right_width_0_height_0_subtile_19__pin_sc_out_0_),
		.ccff_tail(grid_io_left_2_ccff_tail));

	grid_io_left grid_io_left_1__4_ (
		.test_en(test_en),
		.scan_mode(scan_mode),
		.scan_clk(scan_clk),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.CFG_DONE(CFG_DONE),
		.gfpga_pad_QL_PREIO_A2F(gfpga_pad_QL_PREIO_A2F[60:79]),
		.gfpga_pad_QL_PREIO_F2A(gfpga_pad_QL_PREIO_F2A[60:79]),
		.gfpga_pad_QL_PREIO_F2A_DEF0(gfpga_pad_QL_PREIO_F2A_DEF0[60:79]),
		.gfpga_pad_QL_PREIO_F2A_DEF1(gfpga_pad_QL_PREIO_F2A_DEF1[60:79]),
		.gfpga_pad_QL_PREIO_F2A_CLK(gfpga_pad_QL_PREIO_F2A_CLK[60:79]),
		.right_width_0_height_0_subtile_0__pin_f2a_i_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_0__pin_sc_in_0_(grid_io_left_1__4__undriven_right_width_0_height_0_subtile_0__pin_sc_in_0_),
		.right_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_1__pin_f2a_i_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_1__pin_sc_in_0_(grid_io_left_1__4__undriven_right_width_0_height_0_subtile_1__pin_sc_in_0_),
		.right_width_0_height_0_subtile_1__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_1__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_1__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_1__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_1__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_1__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_2__pin_f2a_i_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_2__pin_sc_in_0_(grid_io_left_1__4__undriven_right_width_0_height_0_subtile_2__pin_sc_in_0_),
		.right_width_0_height_0_subtile_2__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_2__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_2__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_2__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_2__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_2__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_3__pin_f2a_i_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_3__pin_sc_in_0_(grid_io_left_1__4__undriven_right_width_0_height_0_subtile_3__pin_sc_in_0_),
		.right_width_0_height_0_subtile_3__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_3__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_3__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_3__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_3__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_3__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_4__pin_f2a_i_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_4__pin_sc_in_0_(grid_io_left_1__4__undriven_right_width_0_height_0_subtile_4__pin_sc_in_0_),
		.right_width_0_height_0_subtile_4__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_4__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_4__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_4__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_4__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_4__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_5__pin_f2a_i_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_5__pin_sc_in_0_(grid_io_left_1__4__undriven_right_width_0_height_0_subtile_5__pin_sc_in_0_),
		.right_width_0_height_0_subtile_5__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_5__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_5__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_5__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_5__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_5__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_6__pin_f2a_i_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_6__pin_sc_in_0_(grid_io_left_1__4__undriven_right_width_0_height_0_subtile_6__pin_sc_in_0_),
		.right_width_0_height_0_subtile_6__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_6__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_6__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_6__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_6__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_6__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_7__pin_f2a_i_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_7__pin_sc_in_0_(grid_io_left_1__4__undriven_right_width_0_height_0_subtile_7__pin_sc_in_0_),
		.right_width_0_height_0_subtile_7__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_7__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_7__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_7__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_7__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_7__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_8__pin_f2a_i_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_8__pin_sc_in_0_(grid_io_left_1__4__undriven_right_width_0_height_0_subtile_8__pin_sc_in_0_),
		.right_width_0_height_0_subtile_8__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_8__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_8__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_8__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_8__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_8__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_9__pin_f2a_i_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_9__pin_sc_in_0_(grid_io_left_1__4__undriven_right_width_0_height_0_subtile_9__pin_sc_in_0_),
		.right_width_0_height_0_subtile_9__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_9__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_9__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_9__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_9__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_9__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_10__pin_f2a_i_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_10__pin_sc_in_0_(grid_io_left_1__4__undriven_right_width_0_height_0_subtile_10__pin_sc_in_0_),
		.right_width_0_height_0_subtile_10__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_10__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_10__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_10__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_10__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_10__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_11__pin_f2a_i_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_11__pin_sc_in_0_(grid_io_left_1__4__undriven_right_width_0_height_0_subtile_11__pin_sc_in_0_),
		.right_width_0_height_0_subtile_11__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_11__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_11__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_11__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_11__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_11__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_12__pin_f2a_i_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_12__pin_sc_in_0_(grid_io_left_1__4__undriven_right_width_0_height_0_subtile_12__pin_sc_in_0_),
		.right_width_0_height_0_subtile_12__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_12__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_12__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_12__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_12__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_12__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_13__pin_f2a_i_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_13__pin_sc_in_0_(grid_io_left_1__4__undriven_right_width_0_height_0_subtile_13__pin_sc_in_0_),
		.right_width_0_height_0_subtile_13__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_13__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_13__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_13__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_13__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_13__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_14__pin_f2a_i_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_14__pin_sc_in_0_(grid_io_left_1__4__undriven_right_width_0_height_0_subtile_14__pin_sc_in_0_),
		.right_width_0_height_0_subtile_14__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_14__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_14__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_14__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_14__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_14__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_15__pin_f2a_i_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_15__pin_sc_in_0_(grid_io_left_1__4__undriven_right_width_0_height_0_subtile_15__pin_sc_in_0_),
		.right_width_0_height_0_subtile_15__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_15__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_15__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_15__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_15__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_15__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_16__pin_f2a_i_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_16__pin_sc_in_0_(grid_io_left_1__4__undriven_right_width_0_height_0_subtile_16__pin_sc_in_0_),
		.right_width_0_height_0_subtile_16__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_16__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_16__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_16__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_16__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_16__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_17__pin_f2a_i_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_17__pin_sc_in_0_(grid_io_left_1__4__undriven_right_width_0_height_0_subtile_17__pin_sc_in_0_),
		.right_width_0_height_0_subtile_17__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_17__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_17__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_17__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_17__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_17__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_18__pin_f2a_i_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_18__pin_sc_in_0_(grid_io_left_1__4__undriven_right_width_0_height_0_subtile_18__pin_sc_in_0_),
		.right_width_0_height_0_subtile_18__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_18__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_18__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_18__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_18__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_18__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_19__pin_f2a_i_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_19__pin_sc_in_0_(grid_io_left_1__4__undriven_right_width_0_height_0_subtile_19__pin_sc_in_0_),
		.right_width_0_height_0_subtile_19__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_19__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_19__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_19__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_19__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_19__pin_clk_3_(clk[3]),
		.ccff_head(cby_1__1__3_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_0__pin_sc_out_0_(grid_io_left_1__4__undriven_right_width_0_height_0_subtile_0__pin_sc_out_0_),
		.right_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_1__pin_sc_out_0_(grid_io_left_1__4__undriven_right_width_0_height_0_subtile_1__pin_sc_out_0_),
		.right_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_2__pin_sc_out_0_(grid_io_left_1__4__undriven_right_width_0_height_0_subtile_2__pin_sc_out_0_),
		.right_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_3__pin_sc_out_0_(grid_io_left_1__4__undriven_right_width_0_height_0_subtile_3__pin_sc_out_0_),
		.right_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_4__pin_sc_out_0_(grid_io_left_1__4__undriven_right_width_0_height_0_subtile_4__pin_sc_out_0_),
		.right_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_5__pin_sc_out_0_(grid_io_left_1__4__undriven_right_width_0_height_0_subtile_5__pin_sc_out_0_),
		.right_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_6__pin_sc_out_0_(grid_io_left_1__4__undriven_right_width_0_height_0_subtile_6__pin_sc_out_0_),
		.right_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_7__pin_sc_out_0_(grid_io_left_1__4__undriven_right_width_0_height_0_subtile_7__pin_sc_out_0_),
		.right_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_8__pin_sc_out_0_(grid_io_left_1__4__undriven_right_width_0_height_0_subtile_8__pin_sc_out_0_),
		.right_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_9__pin_sc_out_0_(grid_io_left_1__4__undriven_right_width_0_height_0_subtile_9__pin_sc_out_0_),
		.right_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_10__pin_sc_out_0_(grid_io_left_1__4__undriven_right_width_0_height_0_subtile_10__pin_sc_out_0_),
		.right_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_11__pin_sc_out_0_(grid_io_left_1__4__undriven_right_width_0_height_0_subtile_11__pin_sc_out_0_),
		.right_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_12__pin_sc_out_0_(grid_io_left_1__4__undriven_right_width_0_height_0_subtile_12__pin_sc_out_0_),
		.right_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_13__pin_sc_out_0_(grid_io_left_1__4__undriven_right_width_0_height_0_subtile_13__pin_sc_out_0_),
		.right_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_14__pin_sc_out_0_(grid_io_left_1__4__undriven_right_width_0_height_0_subtile_14__pin_sc_out_0_),
		.right_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_15__pin_sc_out_0_(grid_io_left_1__4__undriven_right_width_0_height_0_subtile_15__pin_sc_out_0_),
		.right_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_16__pin_sc_out_0_(grid_io_left_1__4__undriven_right_width_0_height_0_subtile_16__pin_sc_out_0_),
		.right_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_17__pin_sc_out_0_(grid_io_left_1__4__undriven_right_width_0_height_0_subtile_17__pin_sc_out_0_),
		.right_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_18__pin_sc_out_0_(grid_io_left_1__4__undriven_right_width_0_height_0_subtile_18__pin_sc_out_0_),
		.right_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_19__pin_sc_out_0_(grid_io_left_1__4__undriven_right_width_0_height_0_subtile_19__pin_sc_out_0_),
		.ccff_tail(grid_io_left_3_ccff_tail));

	grid_io_left grid_io_left_1__5_ (
		.test_en(test_en),
		.scan_mode(scan_mode),
		.scan_clk(scan_clk),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.CFG_DONE(CFG_DONE),
		.gfpga_pad_QL_PREIO_A2F(gfpga_pad_QL_PREIO_A2F[80:99]),
		.gfpga_pad_QL_PREIO_F2A(gfpga_pad_QL_PREIO_F2A[80:99]),
		.gfpga_pad_QL_PREIO_F2A_DEF0(gfpga_pad_QL_PREIO_F2A_DEF0[80:99]),
		.gfpga_pad_QL_PREIO_F2A_DEF1(gfpga_pad_QL_PREIO_F2A_DEF1[80:99]),
		.gfpga_pad_QL_PREIO_F2A_CLK(gfpga_pad_QL_PREIO_F2A_CLK[80:99]),
		.right_width_0_height_0_subtile_0__pin_f2a_i_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_0__pin_sc_in_0_(grid_io_left_1__5__undriven_right_width_0_height_0_subtile_0__pin_sc_in_0_),
		.right_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_1__pin_f2a_i_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_1__pin_sc_in_0_(grid_io_left_1__5__undriven_right_width_0_height_0_subtile_1__pin_sc_in_0_),
		.right_width_0_height_0_subtile_1__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_1__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_1__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_1__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_1__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_1__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_2__pin_f2a_i_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_2__pin_sc_in_0_(grid_io_left_1__5__undriven_right_width_0_height_0_subtile_2__pin_sc_in_0_),
		.right_width_0_height_0_subtile_2__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_2__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_2__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_2__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_2__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_2__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_3__pin_f2a_i_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_3__pin_sc_in_0_(grid_io_left_1__5__undriven_right_width_0_height_0_subtile_3__pin_sc_in_0_),
		.right_width_0_height_0_subtile_3__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_3__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_3__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_3__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_3__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_3__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_4__pin_f2a_i_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_4__pin_sc_in_0_(grid_io_left_1__5__undriven_right_width_0_height_0_subtile_4__pin_sc_in_0_),
		.right_width_0_height_0_subtile_4__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_4__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_4__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_4__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_4__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_4__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_5__pin_f2a_i_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_5__pin_sc_in_0_(grid_io_left_1__5__undriven_right_width_0_height_0_subtile_5__pin_sc_in_0_),
		.right_width_0_height_0_subtile_5__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_5__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_5__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_5__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_5__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_5__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_6__pin_f2a_i_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_6__pin_sc_in_0_(grid_io_left_1__5__undriven_right_width_0_height_0_subtile_6__pin_sc_in_0_),
		.right_width_0_height_0_subtile_6__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_6__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_6__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_6__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_6__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_6__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_7__pin_f2a_i_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_7__pin_sc_in_0_(grid_io_left_1__5__undriven_right_width_0_height_0_subtile_7__pin_sc_in_0_),
		.right_width_0_height_0_subtile_7__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_7__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_7__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_7__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_7__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_7__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_8__pin_f2a_i_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_8__pin_sc_in_0_(grid_io_left_1__5__undriven_right_width_0_height_0_subtile_8__pin_sc_in_0_),
		.right_width_0_height_0_subtile_8__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_8__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_8__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_8__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_8__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_8__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_9__pin_f2a_i_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_9__pin_sc_in_0_(grid_io_left_1__5__undriven_right_width_0_height_0_subtile_9__pin_sc_in_0_),
		.right_width_0_height_0_subtile_9__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_9__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_9__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_9__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_9__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_9__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_10__pin_f2a_i_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_10__pin_sc_in_0_(grid_io_left_1__5__undriven_right_width_0_height_0_subtile_10__pin_sc_in_0_),
		.right_width_0_height_0_subtile_10__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_10__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_10__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_10__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_10__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_10__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_11__pin_f2a_i_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_11__pin_sc_in_0_(grid_io_left_1__5__undriven_right_width_0_height_0_subtile_11__pin_sc_in_0_),
		.right_width_0_height_0_subtile_11__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_11__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_11__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_11__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_11__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_11__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_12__pin_f2a_i_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_12__pin_sc_in_0_(grid_io_left_1__5__undriven_right_width_0_height_0_subtile_12__pin_sc_in_0_),
		.right_width_0_height_0_subtile_12__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_12__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_12__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_12__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_12__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_12__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_13__pin_f2a_i_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_13__pin_sc_in_0_(grid_io_left_1__5__undriven_right_width_0_height_0_subtile_13__pin_sc_in_0_),
		.right_width_0_height_0_subtile_13__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_13__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_13__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_13__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_13__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_13__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_14__pin_f2a_i_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_14__pin_sc_in_0_(grid_io_left_1__5__undriven_right_width_0_height_0_subtile_14__pin_sc_in_0_),
		.right_width_0_height_0_subtile_14__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_14__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_14__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_14__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_14__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_14__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_15__pin_f2a_i_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_15__pin_sc_in_0_(grid_io_left_1__5__undriven_right_width_0_height_0_subtile_15__pin_sc_in_0_),
		.right_width_0_height_0_subtile_15__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_15__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_15__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_15__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_15__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_15__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_16__pin_f2a_i_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_16__pin_sc_in_0_(grid_io_left_1__5__undriven_right_width_0_height_0_subtile_16__pin_sc_in_0_),
		.right_width_0_height_0_subtile_16__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_16__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_16__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_16__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_16__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_16__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_17__pin_f2a_i_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_17__pin_sc_in_0_(grid_io_left_1__5__undriven_right_width_0_height_0_subtile_17__pin_sc_in_0_),
		.right_width_0_height_0_subtile_17__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_17__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_17__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_17__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_17__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_17__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_18__pin_f2a_i_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_18__pin_sc_in_0_(grid_io_left_1__5__undriven_right_width_0_height_0_subtile_18__pin_sc_in_0_),
		.right_width_0_height_0_subtile_18__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_18__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_18__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_18__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_18__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_18__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_19__pin_f2a_i_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_19__pin_sc_in_0_(grid_io_left_1__5__undriven_right_width_0_height_0_subtile_19__pin_sc_in_0_),
		.right_width_0_height_0_subtile_19__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_19__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_19__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_19__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_19__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_19__pin_clk_3_(clk[3]),
		.ccff_head(cby_1__1__4_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_0__pin_sc_out_0_(grid_io_left_1__5__undriven_right_width_0_height_0_subtile_0__pin_sc_out_0_),
		.right_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_1__pin_sc_out_0_(grid_io_left_1__5__undriven_right_width_0_height_0_subtile_1__pin_sc_out_0_),
		.right_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_2__pin_sc_out_0_(grid_io_left_1__5__undriven_right_width_0_height_0_subtile_2__pin_sc_out_0_),
		.right_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_3__pin_sc_out_0_(grid_io_left_1__5__undriven_right_width_0_height_0_subtile_3__pin_sc_out_0_),
		.right_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_4__pin_sc_out_0_(grid_io_left_1__5__undriven_right_width_0_height_0_subtile_4__pin_sc_out_0_),
		.right_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_5__pin_sc_out_0_(grid_io_left_1__5__undriven_right_width_0_height_0_subtile_5__pin_sc_out_0_),
		.right_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_6__pin_sc_out_0_(grid_io_left_1__5__undriven_right_width_0_height_0_subtile_6__pin_sc_out_0_),
		.right_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_7__pin_sc_out_0_(grid_io_left_1__5__undriven_right_width_0_height_0_subtile_7__pin_sc_out_0_),
		.right_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_8__pin_sc_out_0_(grid_io_left_1__5__undriven_right_width_0_height_0_subtile_8__pin_sc_out_0_),
		.right_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_9__pin_sc_out_0_(grid_io_left_1__5__undriven_right_width_0_height_0_subtile_9__pin_sc_out_0_),
		.right_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_10__pin_sc_out_0_(grid_io_left_1__5__undriven_right_width_0_height_0_subtile_10__pin_sc_out_0_),
		.right_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_11__pin_sc_out_0_(grid_io_left_1__5__undriven_right_width_0_height_0_subtile_11__pin_sc_out_0_),
		.right_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_12__pin_sc_out_0_(grid_io_left_1__5__undriven_right_width_0_height_0_subtile_12__pin_sc_out_0_),
		.right_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_13__pin_sc_out_0_(grid_io_left_1__5__undriven_right_width_0_height_0_subtile_13__pin_sc_out_0_),
		.right_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_14__pin_sc_out_0_(grid_io_left_1__5__undriven_right_width_0_height_0_subtile_14__pin_sc_out_0_),
		.right_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_15__pin_sc_out_0_(grid_io_left_1__5__undriven_right_width_0_height_0_subtile_15__pin_sc_out_0_),
		.right_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_16__pin_sc_out_0_(grid_io_left_1__5__undriven_right_width_0_height_0_subtile_16__pin_sc_out_0_),
		.right_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_17__pin_sc_out_0_(grid_io_left_1__5__undriven_right_width_0_height_0_subtile_17__pin_sc_out_0_),
		.right_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_18__pin_sc_out_0_(grid_io_left_1__5__undriven_right_width_0_height_0_subtile_18__pin_sc_out_0_),
		.right_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_19__pin_sc_out_0_(grid_io_left_1__5__undriven_right_width_0_height_0_subtile_19__pin_sc_out_0_),
		.ccff_tail(grid_io_left_4_ccff_tail));

	grid_io_left grid_io_left_1__6_ (
		.test_en(test_en),
		.scan_mode(scan_mode),
		.scan_clk(scan_clk),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.CFG_DONE(CFG_DONE),
		.gfpga_pad_QL_PREIO_A2F(gfpga_pad_QL_PREIO_A2F[100:119]),
		.gfpga_pad_QL_PREIO_F2A(gfpga_pad_QL_PREIO_F2A[100:119]),
		.gfpga_pad_QL_PREIO_F2A_DEF0(gfpga_pad_QL_PREIO_F2A_DEF0[100:119]),
		.gfpga_pad_QL_PREIO_F2A_DEF1(gfpga_pad_QL_PREIO_F2A_DEF1[100:119]),
		.gfpga_pad_QL_PREIO_F2A_CLK(gfpga_pad_QL_PREIO_F2A_CLK[100:119]),
		.right_width_0_height_0_subtile_0__pin_f2a_i_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_0__pin_sc_in_0_(grid_io_left_1__6__undriven_right_width_0_height_0_subtile_0__pin_sc_in_0_),
		.right_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_1__pin_f2a_i_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_1__pin_sc_in_0_(grid_io_left_1__6__undriven_right_width_0_height_0_subtile_1__pin_sc_in_0_),
		.right_width_0_height_0_subtile_1__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_1__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_1__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_1__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_1__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_1__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_2__pin_f2a_i_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_2__pin_sc_in_0_(grid_io_left_1__6__undriven_right_width_0_height_0_subtile_2__pin_sc_in_0_),
		.right_width_0_height_0_subtile_2__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_2__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_2__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_2__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_2__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_2__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_3__pin_f2a_i_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_3__pin_sc_in_0_(grid_io_left_1__6__undriven_right_width_0_height_0_subtile_3__pin_sc_in_0_),
		.right_width_0_height_0_subtile_3__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_3__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_3__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_3__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_3__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_3__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_4__pin_f2a_i_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_4__pin_sc_in_0_(grid_io_left_1__6__undriven_right_width_0_height_0_subtile_4__pin_sc_in_0_),
		.right_width_0_height_0_subtile_4__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_4__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_4__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_4__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_4__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_4__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_5__pin_f2a_i_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_5__pin_sc_in_0_(grid_io_left_1__6__undriven_right_width_0_height_0_subtile_5__pin_sc_in_0_),
		.right_width_0_height_0_subtile_5__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_5__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_5__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_5__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_5__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_5__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_6__pin_f2a_i_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_6__pin_sc_in_0_(grid_io_left_1__6__undriven_right_width_0_height_0_subtile_6__pin_sc_in_0_),
		.right_width_0_height_0_subtile_6__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_6__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_6__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_6__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_6__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_6__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_7__pin_f2a_i_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_7__pin_sc_in_0_(grid_io_left_1__6__undriven_right_width_0_height_0_subtile_7__pin_sc_in_0_),
		.right_width_0_height_0_subtile_7__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_7__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_7__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_7__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_7__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_7__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_8__pin_f2a_i_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_8__pin_sc_in_0_(grid_io_left_1__6__undriven_right_width_0_height_0_subtile_8__pin_sc_in_0_),
		.right_width_0_height_0_subtile_8__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_8__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_8__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_8__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_8__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_8__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_9__pin_f2a_i_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_9__pin_sc_in_0_(grid_io_left_1__6__undriven_right_width_0_height_0_subtile_9__pin_sc_in_0_),
		.right_width_0_height_0_subtile_9__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_9__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_9__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_9__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_9__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_9__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_10__pin_f2a_i_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_10__pin_sc_in_0_(grid_io_left_1__6__undriven_right_width_0_height_0_subtile_10__pin_sc_in_0_),
		.right_width_0_height_0_subtile_10__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_10__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_10__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_10__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_10__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_10__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_11__pin_f2a_i_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_11__pin_sc_in_0_(grid_io_left_1__6__undriven_right_width_0_height_0_subtile_11__pin_sc_in_0_),
		.right_width_0_height_0_subtile_11__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_11__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_11__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_11__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_11__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_11__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_12__pin_f2a_i_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_12__pin_sc_in_0_(grid_io_left_1__6__undriven_right_width_0_height_0_subtile_12__pin_sc_in_0_),
		.right_width_0_height_0_subtile_12__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_12__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_12__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_12__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_12__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_12__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_13__pin_f2a_i_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_13__pin_sc_in_0_(grid_io_left_1__6__undriven_right_width_0_height_0_subtile_13__pin_sc_in_0_),
		.right_width_0_height_0_subtile_13__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_13__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_13__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_13__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_13__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_13__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_14__pin_f2a_i_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_14__pin_sc_in_0_(grid_io_left_1__6__undriven_right_width_0_height_0_subtile_14__pin_sc_in_0_),
		.right_width_0_height_0_subtile_14__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_14__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_14__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_14__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_14__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_14__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_15__pin_f2a_i_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_15__pin_sc_in_0_(grid_io_left_1__6__undriven_right_width_0_height_0_subtile_15__pin_sc_in_0_),
		.right_width_0_height_0_subtile_15__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_15__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_15__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_15__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_15__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_15__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_16__pin_f2a_i_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_16__pin_sc_in_0_(grid_io_left_1__6__undriven_right_width_0_height_0_subtile_16__pin_sc_in_0_),
		.right_width_0_height_0_subtile_16__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_16__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_16__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_16__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_16__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_16__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_17__pin_f2a_i_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_17__pin_sc_in_0_(grid_io_left_1__6__undriven_right_width_0_height_0_subtile_17__pin_sc_in_0_),
		.right_width_0_height_0_subtile_17__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_17__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_17__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_17__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_17__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_17__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_18__pin_f2a_i_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_18__pin_sc_in_0_(grid_io_left_1__6__undriven_right_width_0_height_0_subtile_18__pin_sc_in_0_),
		.right_width_0_height_0_subtile_18__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_18__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_18__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_18__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_18__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_18__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_19__pin_f2a_i_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_19__pin_sc_in_0_(grid_io_left_1__6__undriven_right_width_0_height_0_subtile_19__pin_sc_in_0_),
		.right_width_0_height_0_subtile_19__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_19__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_19__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_19__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_19__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_19__pin_clk_3_(clk[3]),
		.ccff_head(cby_1__1__5_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_0__pin_sc_out_0_(grid_io_left_1__6__undriven_right_width_0_height_0_subtile_0__pin_sc_out_0_),
		.right_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_1__pin_sc_out_0_(grid_io_left_1__6__undriven_right_width_0_height_0_subtile_1__pin_sc_out_0_),
		.right_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_2__pin_sc_out_0_(grid_io_left_1__6__undriven_right_width_0_height_0_subtile_2__pin_sc_out_0_),
		.right_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_3__pin_sc_out_0_(grid_io_left_1__6__undriven_right_width_0_height_0_subtile_3__pin_sc_out_0_),
		.right_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_4__pin_sc_out_0_(grid_io_left_1__6__undriven_right_width_0_height_0_subtile_4__pin_sc_out_0_),
		.right_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_5__pin_sc_out_0_(grid_io_left_1__6__undriven_right_width_0_height_0_subtile_5__pin_sc_out_0_),
		.right_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_6__pin_sc_out_0_(grid_io_left_1__6__undriven_right_width_0_height_0_subtile_6__pin_sc_out_0_),
		.right_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_7__pin_sc_out_0_(grid_io_left_1__6__undriven_right_width_0_height_0_subtile_7__pin_sc_out_0_),
		.right_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_8__pin_sc_out_0_(grid_io_left_1__6__undriven_right_width_0_height_0_subtile_8__pin_sc_out_0_),
		.right_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_9__pin_sc_out_0_(grid_io_left_1__6__undriven_right_width_0_height_0_subtile_9__pin_sc_out_0_),
		.right_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_10__pin_sc_out_0_(grid_io_left_1__6__undriven_right_width_0_height_0_subtile_10__pin_sc_out_0_),
		.right_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_11__pin_sc_out_0_(grid_io_left_1__6__undriven_right_width_0_height_0_subtile_11__pin_sc_out_0_),
		.right_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_12__pin_sc_out_0_(grid_io_left_1__6__undriven_right_width_0_height_0_subtile_12__pin_sc_out_0_),
		.right_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_13__pin_sc_out_0_(grid_io_left_1__6__undriven_right_width_0_height_0_subtile_13__pin_sc_out_0_),
		.right_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_14__pin_sc_out_0_(grid_io_left_1__6__undriven_right_width_0_height_0_subtile_14__pin_sc_out_0_),
		.right_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_15__pin_sc_out_0_(grid_io_left_1__6__undriven_right_width_0_height_0_subtile_15__pin_sc_out_0_),
		.right_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_16__pin_sc_out_0_(grid_io_left_1__6__undriven_right_width_0_height_0_subtile_16__pin_sc_out_0_),
		.right_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_17__pin_sc_out_0_(grid_io_left_1__6__undriven_right_width_0_height_0_subtile_17__pin_sc_out_0_),
		.right_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_18__pin_sc_out_0_(grid_io_left_1__6__undriven_right_width_0_height_0_subtile_18__pin_sc_out_0_),
		.right_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_19__pin_sc_out_0_(grid_io_left_1__6__undriven_right_width_0_height_0_subtile_19__pin_sc_out_0_),
		.ccff_tail(grid_io_left_5_ccff_tail));

	grid_io_left grid_io_left_1__7_ (
		.test_en(test_en),
		.scan_mode(scan_mode),
		.scan_clk(scan_clk),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.CFG_DONE(CFG_DONE),
		.gfpga_pad_QL_PREIO_A2F(gfpga_pad_QL_PREIO_A2F[120:139]),
		.gfpga_pad_QL_PREIO_F2A(gfpga_pad_QL_PREIO_F2A[120:139]),
		.gfpga_pad_QL_PREIO_F2A_DEF0(gfpga_pad_QL_PREIO_F2A_DEF0[120:139]),
		.gfpga_pad_QL_PREIO_F2A_DEF1(gfpga_pad_QL_PREIO_F2A_DEF1[120:139]),
		.gfpga_pad_QL_PREIO_F2A_CLK(gfpga_pad_QL_PREIO_F2A_CLK[120:139]),
		.right_width_0_height_0_subtile_0__pin_f2a_i_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_0__pin_sc_in_0_(grid_io_left_1__7__undriven_right_width_0_height_0_subtile_0__pin_sc_in_0_),
		.right_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_1__pin_f2a_i_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_1__pin_sc_in_0_(grid_io_left_1__7__undriven_right_width_0_height_0_subtile_1__pin_sc_in_0_),
		.right_width_0_height_0_subtile_1__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_1__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_1__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_1__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_1__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_1__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_2__pin_f2a_i_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_2__pin_sc_in_0_(grid_io_left_1__7__undriven_right_width_0_height_0_subtile_2__pin_sc_in_0_),
		.right_width_0_height_0_subtile_2__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_2__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_2__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_2__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_2__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_2__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_3__pin_f2a_i_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_3__pin_sc_in_0_(grid_io_left_1__7__undriven_right_width_0_height_0_subtile_3__pin_sc_in_0_),
		.right_width_0_height_0_subtile_3__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_3__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_3__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_3__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_3__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_3__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_4__pin_f2a_i_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_4__pin_sc_in_0_(grid_io_left_1__7__undriven_right_width_0_height_0_subtile_4__pin_sc_in_0_),
		.right_width_0_height_0_subtile_4__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_4__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_4__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_4__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_4__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_4__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_5__pin_f2a_i_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_5__pin_sc_in_0_(grid_io_left_1__7__undriven_right_width_0_height_0_subtile_5__pin_sc_in_0_),
		.right_width_0_height_0_subtile_5__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_5__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_5__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_5__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_5__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_5__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_6__pin_f2a_i_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_6__pin_sc_in_0_(grid_io_left_1__7__undriven_right_width_0_height_0_subtile_6__pin_sc_in_0_),
		.right_width_0_height_0_subtile_6__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_6__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_6__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_6__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_6__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_6__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_7__pin_f2a_i_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_7__pin_sc_in_0_(grid_io_left_1__7__undriven_right_width_0_height_0_subtile_7__pin_sc_in_0_),
		.right_width_0_height_0_subtile_7__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_7__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_7__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_7__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_7__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_7__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_8__pin_f2a_i_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_8__pin_sc_in_0_(grid_io_left_1__7__undriven_right_width_0_height_0_subtile_8__pin_sc_in_0_),
		.right_width_0_height_0_subtile_8__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_8__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_8__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_8__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_8__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_8__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_9__pin_f2a_i_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_9__pin_sc_in_0_(grid_io_left_1__7__undriven_right_width_0_height_0_subtile_9__pin_sc_in_0_),
		.right_width_0_height_0_subtile_9__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_9__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_9__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_9__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_9__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_9__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_10__pin_f2a_i_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_10__pin_sc_in_0_(grid_io_left_1__7__undriven_right_width_0_height_0_subtile_10__pin_sc_in_0_),
		.right_width_0_height_0_subtile_10__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_10__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_10__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_10__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_10__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_10__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_11__pin_f2a_i_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_11__pin_sc_in_0_(grid_io_left_1__7__undriven_right_width_0_height_0_subtile_11__pin_sc_in_0_),
		.right_width_0_height_0_subtile_11__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_11__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_11__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_11__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_11__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_11__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_12__pin_f2a_i_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_12__pin_sc_in_0_(grid_io_left_1__7__undriven_right_width_0_height_0_subtile_12__pin_sc_in_0_),
		.right_width_0_height_0_subtile_12__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_12__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_12__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_12__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_12__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_12__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_13__pin_f2a_i_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_13__pin_sc_in_0_(grid_io_left_1__7__undriven_right_width_0_height_0_subtile_13__pin_sc_in_0_),
		.right_width_0_height_0_subtile_13__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_13__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_13__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_13__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_13__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_13__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_14__pin_f2a_i_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_14__pin_sc_in_0_(grid_io_left_1__7__undriven_right_width_0_height_0_subtile_14__pin_sc_in_0_),
		.right_width_0_height_0_subtile_14__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_14__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_14__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_14__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_14__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_14__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_15__pin_f2a_i_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_15__pin_sc_in_0_(grid_io_left_1__7__undriven_right_width_0_height_0_subtile_15__pin_sc_in_0_),
		.right_width_0_height_0_subtile_15__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_15__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_15__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_15__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_15__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_15__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_16__pin_f2a_i_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_16__pin_sc_in_0_(grid_io_left_1__7__undriven_right_width_0_height_0_subtile_16__pin_sc_in_0_),
		.right_width_0_height_0_subtile_16__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_16__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_16__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_16__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_16__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_16__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_17__pin_f2a_i_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_17__pin_sc_in_0_(grid_io_left_1__7__undriven_right_width_0_height_0_subtile_17__pin_sc_in_0_),
		.right_width_0_height_0_subtile_17__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_17__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_17__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_17__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_17__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_17__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_18__pin_f2a_i_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_18__pin_sc_in_0_(grid_io_left_1__7__undriven_right_width_0_height_0_subtile_18__pin_sc_in_0_),
		.right_width_0_height_0_subtile_18__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_18__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_18__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_18__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_18__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_18__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_19__pin_f2a_i_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_19__pin_sc_in_0_(grid_io_left_1__7__undriven_right_width_0_height_0_subtile_19__pin_sc_in_0_),
		.right_width_0_height_0_subtile_19__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_19__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_19__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_19__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_19__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_19__pin_clk_3_(clk[3]),
		.ccff_head(cby_1__1__6_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_0__pin_sc_out_0_(grid_io_left_1__7__undriven_right_width_0_height_0_subtile_0__pin_sc_out_0_),
		.right_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_1__pin_sc_out_0_(grid_io_left_1__7__undriven_right_width_0_height_0_subtile_1__pin_sc_out_0_),
		.right_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_2__pin_sc_out_0_(grid_io_left_1__7__undriven_right_width_0_height_0_subtile_2__pin_sc_out_0_),
		.right_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_3__pin_sc_out_0_(grid_io_left_1__7__undriven_right_width_0_height_0_subtile_3__pin_sc_out_0_),
		.right_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_4__pin_sc_out_0_(grid_io_left_1__7__undriven_right_width_0_height_0_subtile_4__pin_sc_out_0_),
		.right_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_5__pin_sc_out_0_(grid_io_left_1__7__undriven_right_width_0_height_0_subtile_5__pin_sc_out_0_),
		.right_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_6__pin_sc_out_0_(grid_io_left_1__7__undriven_right_width_0_height_0_subtile_6__pin_sc_out_0_),
		.right_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_7__pin_sc_out_0_(grid_io_left_1__7__undriven_right_width_0_height_0_subtile_7__pin_sc_out_0_),
		.right_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_8__pin_sc_out_0_(grid_io_left_1__7__undriven_right_width_0_height_0_subtile_8__pin_sc_out_0_),
		.right_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_9__pin_sc_out_0_(grid_io_left_1__7__undriven_right_width_0_height_0_subtile_9__pin_sc_out_0_),
		.right_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_10__pin_sc_out_0_(grid_io_left_1__7__undriven_right_width_0_height_0_subtile_10__pin_sc_out_0_),
		.right_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_11__pin_sc_out_0_(grid_io_left_1__7__undriven_right_width_0_height_0_subtile_11__pin_sc_out_0_),
		.right_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_12__pin_sc_out_0_(grid_io_left_1__7__undriven_right_width_0_height_0_subtile_12__pin_sc_out_0_),
		.right_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_13__pin_sc_out_0_(grid_io_left_1__7__undriven_right_width_0_height_0_subtile_13__pin_sc_out_0_),
		.right_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_14__pin_sc_out_0_(grid_io_left_1__7__undriven_right_width_0_height_0_subtile_14__pin_sc_out_0_),
		.right_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_15__pin_sc_out_0_(grid_io_left_1__7__undriven_right_width_0_height_0_subtile_15__pin_sc_out_0_),
		.right_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_16__pin_sc_out_0_(grid_io_left_1__7__undriven_right_width_0_height_0_subtile_16__pin_sc_out_0_),
		.right_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_17__pin_sc_out_0_(grid_io_left_1__7__undriven_right_width_0_height_0_subtile_17__pin_sc_out_0_),
		.right_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_18__pin_sc_out_0_(grid_io_left_1__7__undriven_right_width_0_height_0_subtile_18__pin_sc_out_0_),
		.right_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_19__pin_sc_out_0_(grid_io_left_1__7__undriven_right_width_0_height_0_subtile_19__pin_sc_out_0_),
		.ccff_tail(grid_io_left_6_ccff_tail));

	grid_io_left grid_io_left_1__8_ (
		.test_en(test_en),
		.scan_mode(scan_mode),
		.scan_clk(scan_clk),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.CFG_DONE(CFG_DONE),
		.gfpga_pad_QL_PREIO_A2F(gfpga_pad_QL_PREIO_A2F[140:159]),
		.gfpga_pad_QL_PREIO_F2A(gfpga_pad_QL_PREIO_F2A[140:159]),
		.gfpga_pad_QL_PREIO_F2A_DEF0(gfpga_pad_QL_PREIO_F2A_DEF0[140:159]),
		.gfpga_pad_QL_PREIO_F2A_DEF1(gfpga_pad_QL_PREIO_F2A_DEF1[140:159]),
		.gfpga_pad_QL_PREIO_F2A_CLK(gfpga_pad_QL_PREIO_F2A_CLK[140:159]),
		.right_width_0_height_0_subtile_0__pin_f2a_i_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_0__pin_sc_in_0_(grid_io_left_1__8__undriven_right_width_0_height_0_subtile_0__pin_sc_in_0_),
		.right_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_1__pin_f2a_i_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_1__pin_sc_in_0_(grid_io_left_1__8__undriven_right_width_0_height_0_subtile_1__pin_sc_in_0_),
		.right_width_0_height_0_subtile_1__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_1__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_1__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_1__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_1__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_1__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_2__pin_f2a_i_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_2__pin_sc_in_0_(grid_io_left_1__8__undriven_right_width_0_height_0_subtile_2__pin_sc_in_0_),
		.right_width_0_height_0_subtile_2__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_2__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_2__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_2__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_2__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_2__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_3__pin_f2a_i_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_3__pin_sc_in_0_(grid_io_left_1__8__undriven_right_width_0_height_0_subtile_3__pin_sc_in_0_),
		.right_width_0_height_0_subtile_3__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_3__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_3__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_3__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_3__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_3__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_4__pin_f2a_i_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_4__pin_sc_in_0_(grid_io_left_1__8__undriven_right_width_0_height_0_subtile_4__pin_sc_in_0_),
		.right_width_0_height_0_subtile_4__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_4__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_4__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_4__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_4__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_4__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_5__pin_f2a_i_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_5__pin_sc_in_0_(grid_io_left_1__8__undriven_right_width_0_height_0_subtile_5__pin_sc_in_0_),
		.right_width_0_height_0_subtile_5__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_5__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_5__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_5__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_5__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_5__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_6__pin_f2a_i_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_6__pin_sc_in_0_(grid_io_left_1__8__undriven_right_width_0_height_0_subtile_6__pin_sc_in_0_),
		.right_width_0_height_0_subtile_6__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_6__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_6__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_6__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_6__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_6__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_7__pin_f2a_i_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_7__pin_sc_in_0_(grid_io_left_1__8__undriven_right_width_0_height_0_subtile_7__pin_sc_in_0_),
		.right_width_0_height_0_subtile_7__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_7__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_7__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_7__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_7__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_7__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_8__pin_f2a_i_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_8__pin_sc_in_0_(grid_io_left_1__8__undriven_right_width_0_height_0_subtile_8__pin_sc_in_0_),
		.right_width_0_height_0_subtile_8__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_8__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_8__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_8__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_8__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_8__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_9__pin_f2a_i_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_9__pin_sc_in_0_(grid_io_left_1__8__undriven_right_width_0_height_0_subtile_9__pin_sc_in_0_),
		.right_width_0_height_0_subtile_9__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_9__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_9__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_9__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_9__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_9__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_10__pin_f2a_i_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_10__pin_sc_in_0_(grid_io_left_1__8__undriven_right_width_0_height_0_subtile_10__pin_sc_in_0_),
		.right_width_0_height_0_subtile_10__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_10__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_10__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_10__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_10__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_10__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_11__pin_f2a_i_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_11__pin_sc_in_0_(grid_io_left_1__8__undriven_right_width_0_height_0_subtile_11__pin_sc_in_0_),
		.right_width_0_height_0_subtile_11__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_11__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_11__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_11__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_11__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_11__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_12__pin_f2a_i_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_12__pin_sc_in_0_(grid_io_left_1__8__undriven_right_width_0_height_0_subtile_12__pin_sc_in_0_),
		.right_width_0_height_0_subtile_12__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_12__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_12__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_12__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_12__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_12__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_13__pin_f2a_i_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_13__pin_sc_in_0_(grid_io_left_1__8__undriven_right_width_0_height_0_subtile_13__pin_sc_in_0_),
		.right_width_0_height_0_subtile_13__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_13__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_13__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_13__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_13__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_13__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_14__pin_f2a_i_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_14__pin_sc_in_0_(grid_io_left_1__8__undriven_right_width_0_height_0_subtile_14__pin_sc_in_0_),
		.right_width_0_height_0_subtile_14__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_14__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_14__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_14__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_14__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_14__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_15__pin_f2a_i_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_15__pin_sc_in_0_(grid_io_left_1__8__undriven_right_width_0_height_0_subtile_15__pin_sc_in_0_),
		.right_width_0_height_0_subtile_15__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_15__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_15__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_15__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_15__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_15__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_16__pin_f2a_i_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_16__pin_sc_in_0_(grid_io_left_1__8__undriven_right_width_0_height_0_subtile_16__pin_sc_in_0_),
		.right_width_0_height_0_subtile_16__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_16__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_16__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_16__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_16__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_16__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_17__pin_f2a_i_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_17__pin_sc_in_0_(grid_io_left_1__8__undriven_right_width_0_height_0_subtile_17__pin_sc_in_0_),
		.right_width_0_height_0_subtile_17__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_17__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_17__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_17__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_17__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_17__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_18__pin_f2a_i_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_18__pin_sc_in_0_(grid_io_left_1__8__undriven_right_width_0_height_0_subtile_18__pin_sc_in_0_),
		.right_width_0_height_0_subtile_18__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_18__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_18__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_18__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_18__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_18__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_19__pin_f2a_i_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.right_width_0_height_0_subtile_19__pin_sc_in_0_(grid_io_left_1__8__undriven_right_width_0_height_0_subtile_19__pin_sc_in_0_),
		.right_width_0_height_0_subtile_19__pin_global_reset_0_(global_reset),
		.right_width_0_height_0_subtile_19__pin_scan_reset_0_(scan_reset),
		.right_width_0_height_0_subtile_19__pin_clk_0_(clk[0]),
		.right_width_0_height_0_subtile_19__pin_clk_1_(clk[1]),
		.right_width_0_height_0_subtile_19__pin_clk_2_(clk[2]),
		.right_width_0_height_0_subtile_19__pin_clk_3_(clk[3]),
		.ccff_head(cby_1__1__7_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_0__pin_sc_out_0_(grid_io_left_1__8__undriven_right_width_0_height_0_subtile_0__pin_sc_out_0_),
		.right_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_1__pin_sc_out_0_(grid_io_left_1__8__undriven_right_width_0_height_0_subtile_1__pin_sc_out_0_),
		.right_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_2__pin_sc_out_0_(grid_io_left_1__8__undriven_right_width_0_height_0_subtile_2__pin_sc_out_0_),
		.right_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_3__pin_sc_out_0_(grid_io_left_1__8__undriven_right_width_0_height_0_subtile_3__pin_sc_out_0_),
		.right_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_4__pin_sc_out_0_(grid_io_left_1__8__undriven_right_width_0_height_0_subtile_4__pin_sc_out_0_),
		.right_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_5__pin_sc_out_0_(grid_io_left_1__8__undriven_right_width_0_height_0_subtile_5__pin_sc_out_0_),
		.right_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_6__pin_sc_out_0_(grid_io_left_1__8__undriven_right_width_0_height_0_subtile_6__pin_sc_out_0_),
		.right_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_7__pin_sc_out_0_(grid_io_left_1__8__undriven_right_width_0_height_0_subtile_7__pin_sc_out_0_),
		.right_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_8__pin_sc_out_0_(grid_io_left_1__8__undriven_right_width_0_height_0_subtile_8__pin_sc_out_0_),
		.right_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_9__pin_sc_out_0_(grid_io_left_1__8__undriven_right_width_0_height_0_subtile_9__pin_sc_out_0_),
		.right_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_10__pin_sc_out_0_(grid_io_left_1__8__undriven_right_width_0_height_0_subtile_10__pin_sc_out_0_),
		.right_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_11__pin_sc_out_0_(grid_io_left_1__8__undriven_right_width_0_height_0_subtile_11__pin_sc_out_0_),
		.right_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_12__pin_sc_out_0_(grid_io_left_1__8__undriven_right_width_0_height_0_subtile_12__pin_sc_out_0_),
		.right_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_13__pin_sc_out_0_(grid_io_left_1__8__undriven_right_width_0_height_0_subtile_13__pin_sc_out_0_),
		.right_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_14__pin_sc_out_0_(grid_io_left_1__8__undriven_right_width_0_height_0_subtile_14__pin_sc_out_0_),
		.right_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_15__pin_sc_out_0_(grid_io_left_1__8__undriven_right_width_0_height_0_subtile_15__pin_sc_out_0_),
		.right_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_16__pin_sc_out_0_(grid_io_left_1__8__undriven_right_width_0_height_0_subtile_16__pin_sc_out_0_),
		.right_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_17__pin_sc_out_0_(grid_io_left_1__8__undriven_right_width_0_height_0_subtile_17__pin_sc_out_0_),
		.right_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_18__pin_sc_out_0_(grid_io_left_1__8__undriven_right_width_0_height_0_subtile_18__pin_sc_out_0_),
		.right_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.right_width_0_height_0_subtile_19__pin_sc_out_0_(grid_io_left_1__8__undriven_right_width_0_height_0_subtile_19__pin_sc_out_0_),
		.ccff_tail(ccff_tail[9]));

	grid_io_bottom grid_io_bottom_2__1_ (
		.test_en(test_en),
		.scan_mode(scan_mode),
		.scan_clk(scan_clk),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.CFG_DONE(CFG_DONE),
		.gfpga_pad_QL_PREIO_A2F(gfpga_pad_QL_PREIO_A2F[620:639]),
		.gfpga_pad_QL_PREIO_F2A(gfpga_pad_QL_PREIO_F2A[620:639]),
		.gfpga_pad_QL_PREIO_F2A_DEF0(gfpga_pad_QL_PREIO_F2A_DEF0[620:639]),
		.gfpga_pad_QL_PREIO_F2A_DEF1(gfpga_pad_QL_PREIO_F2A_DEF1[620:639]),
		.gfpga_pad_QL_PREIO_F2A_CLK(gfpga_pad_QL_PREIO_F2A_CLK[620:639]),
		.top_width_0_height_0_subtile_0__pin_f2a_i_0_(cbx_2__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_io_bottom_2__1__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
		.top_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_1__pin_f2a_i_0_(cbx_2__1__0_bottom_grid_top_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_1__pin_sc_in_0_(grid_io_bottom_2__1__undriven_top_width_0_height_0_subtile_1__pin_sc_in_0_),
		.top_width_0_height_0_subtile_1__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_1__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_1__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_1__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_1__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_1__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_2__pin_f2a_i_0_(cbx_2__1__0_bottom_grid_top_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_2__pin_sc_in_0_(grid_io_bottom_2__1__undriven_top_width_0_height_0_subtile_2__pin_sc_in_0_),
		.top_width_0_height_0_subtile_2__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_2__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_2__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_2__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_2__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_2__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_3__pin_f2a_i_0_(cbx_2__1__0_bottom_grid_top_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_3__pin_sc_in_0_(grid_io_bottom_2__1__undriven_top_width_0_height_0_subtile_3__pin_sc_in_0_),
		.top_width_0_height_0_subtile_3__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_3__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_3__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_3__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_3__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_3__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_4__pin_f2a_i_0_(cbx_2__1__0_bottom_grid_top_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_4__pin_sc_in_0_(grid_io_bottom_2__1__undriven_top_width_0_height_0_subtile_4__pin_sc_in_0_),
		.top_width_0_height_0_subtile_4__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_4__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_4__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_4__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_4__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_4__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_5__pin_f2a_i_0_(cbx_2__1__0_bottom_grid_top_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_5__pin_sc_in_0_(grid_io_bottom_2__1__undriven_top_width_0_height_0_subtile_5__pin_sc_in_0_),
		.top_width_0_height_0_subtile_5__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_5__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_5__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_5__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_5__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_5__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_6__pin_f2a_i_0_(cbx_2__1__0_bottom_grid_top_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_6__pin_sc_in_0_(grid_io_bottom_2__1__undriven_top_width_0_height_0_subtile_6__pin_sc_in_0_),
		.top_width_0_height_0_subtile_6__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_6__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_6__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_6__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_6__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_6__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_7__pin_f2a_i_0_(cbx_2__1__0_bottom_grid_top_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_7__pin_sc_in_0_(grid_io_bottom_2__1__undriven_top_width_0_height_0_subtile_7__pin_sc_in_0_),
		.top_width_0_height_0_subtile_7__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_7__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_7__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_7__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_7__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_7__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_8__pin_f2a_i_0_(cbx_2__1__0_bottom_grid_top_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_8__pin_sc_in_0_(grid_io_bottom_2__1__undriven_top_width_0_height_0_subtile_8__pin_sc_in_0_),
		.top_width_0_height_0_subtile_8__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_8__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_8__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_8__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_8__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_8__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_9__pin_f2a_i_0_(cbx_2__1__0_bottom_grid_top_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_9__pin_sc_in_0_(grid_io_bottom_2__1__undriven_top_width_0_height_0_subtile_9__pin_sc_in_0_),
		.top_width_0_height_0_subtile_9__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_9__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_9__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_9__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_9__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_9__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_10__pin_f2a_i_0_(cbx_2__1__0_bottom_grid_top_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_10__pin_sc_in_0_(grid_io_bottom_2__1__undriven_top_width_0_height_0_subtile_10__pin_sc_in_0_),
		.top_width_0_height_0_subtile_10__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_10__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_10__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_10__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_10__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_10__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_11__pin_f2a_i_0_(cbx_2__1__0_bottom_grid_top_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_11__pin_sc_in_0_(grid_io_bottom_2__1__undriven_top_width_0_height_0_subtile_11__pin_sc_in_0_),
		.top_width_0_height_0_subtile_11__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_11__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_11__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_11__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_11__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_11__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_12__pin_f2a_i_0_(cbx_2__1__0_bottom_grid_top_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_12__pin_sc_in_0_(grid_io_bottom_2__1__undriven_top_width_0_height_0_subtile_12__pin_sc_in_0_),
		.top_width_0_height_0_subtile_12__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_12__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_12__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_12__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_12__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_12__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_13__pin_f2a_i_0_(cbx_2__1__0_bottom_grid_top_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_13__pin_sc_in_0_(grid_io_bottom_2__1__undriven_top_width_0_height_0_subtile_13__pin_sc_in_0_),
		.top_width_0_height_0_subtile_13__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_13__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_13__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_13__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_13__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_13__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_14__pin_f2a_i_0_(cbx_2__1__0_bottom_grid_top_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_14__pin_sc_in_0_(grid_io_bottom_2__1__undriven_top_width_0_height_0_subtile_14__pin_sc_in_0_),
		.top_width_0_height_0_subtile_14__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_14__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_14__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_14__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_14__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_14__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_15__pin_f2a_i_0_(cbx_2__1__0_bottom_grid_top_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_15__pin_sc_in_0_(grid_io_bottom_2__1__undriven_top_width_0_height_0_subtile_15__pin_sc_in_0_),
		.top_width_0_height_0_subtile_15__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_15__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_15__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_15__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_15__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_15__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_16__pin_f2a_i_0_(cbx_2__1__0_bottom_grid_top_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_16__pin_sc_in_0_(grid_io_bottom_2__1__undriven_top_width_0_height_0_subtile_16__pin_sc_in_0_),
		.top_width_0_height_0_subtile_16__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_16__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_16__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_16__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_16__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_16__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_17__pin_f2a_i_0_(cbx_2__1__0_bottom_grid_top_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_17__pin_sc_in_0_(grid_io_bottom_2__1__undriven_top_width_0_height_0_subtile_17__pin_sc_in_0_),
		.top_width_0_height_0_subtile_17__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_17__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_17__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_17__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_17__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_17__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_18__pin_f2a_i_0_(cbx_2__1__0_bottom_grid_top_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_18__pin_sc_in_0_(grid_io_bottom_2__1__undriven_top_width_0_height_0_subtile_18__pin_sc_in_0_),
		.top_width_0_height_0_subtile_18__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_18__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_18__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_18__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_18__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_18__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_19__pin_f2a_i_0_(cbx_2__1__0_bottom_grid_top_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_19__pin_sc_in_0_(grid_io_bottom_2__1__undriven_top_width_0_height_0_subtile_19__pin_sc_in_0_),
		.top_width_0_height_0_subtile_19__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_19__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_19__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_19__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_19__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_19__pin_clk_3_(clk[3]),
		.ccff_head(sb_2__0__0_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_0__pin_sc_out_0_(grid_io_bottom_2__1__undriven_top_width_0_height_0_subtile_0__pin_sc_out_0_),
		.top_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_1__pin_sc_out_0_(grid_io_bottom_2__1__undriven_top_width_0_height_0_subtile_1__pin_sc_out_0_),
		.top_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_2__pin_sc_out_0_(grid_io_bottom_2__1__undriven_top_width_0_height_0_subtile_2__pin_sc_out_0_),
		.top_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_3__pin_sc_out_0_(grid_io_bottom_2__1__undriven_top_width_0_height_0_subtile_3__pin_sc_out_0_),
		.top_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_4__pin_sc_out_0_(grid_io_bottom_2__1__undriven_top_width_0_height_0_subtile_4__pin_sc_out_0_),
		.top_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_5__pin_sc_out_0_(grid_io_bottom_2__1__undriven_top_width_0_height_0_subtile_5__pin_sc_out_0_),
		.top_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_6__pin_sc_out_0_(grid_io_bottom_2__1__undriven_top_width_0_height_0_subtile_6__pin_sc_out_0_),
		.top_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_7__pin_sc_out_0_(grid_io_bottom_2__1__undriven_top_width_0_height_0_subtile_7__pin_sc_out_0_),
		.top_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_8__pin_sc_out_0_(grid_io_bottom_2__1__undriven_top_width_0_height_0_subtile_8__pin_sc_out_0_),
		.top_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_9__pin_sc_out_0_(grid_io_bottom_2__1__undriven_top_width_0_height_0_subtile_9__pin_sc_out_0_),
		.top_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_10__pin_sc_out_0_(grid_io_bottom_2__1__undriven_top_width_0_height_0_subtile_10__pin_sc_out_0_),
		.top_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_11__pin_sc_out_0_(grid_io_bottom_2__1__undriven_top_width_0_height_0_subtile_11__pin_sc_out_0_),
		.top_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_12__pin_sc_out_0_(grid_io_bottom_2__1__undriven_top_width_0_height_0_subtile_12__pin_sc_out_0_),
		.top_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_13__pin_sc_out_0_(grid_io_bottom_2__1__undriven_top_width_0_height_0_subtile_13__pin_sc_out_0_),
		.top_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_14__pin_sc_out_0_(grid_io_bottom_2__1__undriven_top_width_0_height_0_subtile_14__pin_sc_out_0_),
		.top_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_15__pin_sc_out_0_(grid_io_bottom_2__1__undriven_top_width_0_height_0_subtile_15__pin_sc_out_0_),
		.top_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_16__pin_sc_out_0_(grid_io_bottom_2__1__undriven_top_width_0_height_0_subtile_16__pin_sc_out_0_),
		.top_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_17__pin_sc_out_0_(grid_io_bottom_2__1__undriven_top_width_0_height_0_subtile_17__pin_sc_out_0_),
		.top_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_18__pin_sc_out_0_(grid_io_bottom_2__1__undriven_top_width_0_height_0_subtile_18__pin_sc_out_0_),
		.top_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_19__pin_sc_out_0_(grid_io_bottom_2__1__undriven_top_width_0_height_0_subtile_19__pin_sc_out_0_),
		.ccff_tail(grid_io_bottom_0_ccff_tail));

	grid_io_bottom grid_io_bottom_3__1_ (
		.test_en(test_en),
		.scan_mode(scan_mode),
		.scan_clk(scan_clk),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.CFG_DONE(CFG_DONE),
		.gfpga_pad_QL_PREIO_A2F(gfpga_pad_QL_PREIO_A2F[600:619]),
		.gfpga_pad_QL_PREIO_F2A(gfpga_pad_QL_PREIO_F2A[600:619]),
		.gfpga_pad_QL_PREIO_F2A_DEF0(gfpga_pad_QL_PREIO_F2A_DEF0[600:619]),
		.gfpga_pad_QL_PREIO_F2A_DEF1(gfpga_pad_QL_PREIO_F2A_DEF1[600:619]),
		.gfpga_pad_QL_PREIO_F2A_CLK(gfpga_pad_QL_PREIO_F2A_CLK[600:619]),
		.top_width_0_height_0_subtile_0__pin_f2a_i_0_(cbx_2__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_io_bottom_3__1__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
		.top_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_1__pin_f2a_i_0_(cbx_2__1__1_bottom_grid_top_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_1__pin_sc_in_0_(grid_io_bottom_3__1__undriven_top_width_0_height_0_subtile_1__pin_sc_in_0_),
		.top_width_0_height_0_subtile_1__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_1__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_1__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_1__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_1__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_1__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_2__pin_f2a_i_0_(cbx_2__1__1_bottom_grid_top_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_2__pin_sc_in_0_(grid_io_bottom_3__1__undriven_top_width_0_height_0_subtile_2__pin_sc_in_0_),
		.top_width_0_height_0_subtile_2__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_2__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_2__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_2__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_2__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_2__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_3__pin_f2a_i_0_(cbx_2__1__1_bottom_grid_top_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_3__pin_sc_in_0_(grid_io_bottom_3__1__undriven_top_width_0_height_0_subtile_3__pin_sc_in_0_),
		.top_width_0_height_0_subtile_3__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_3__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_3__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_3__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_3__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_3__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_4__pin_f2a_i_0_(cbx_2__1__1_bottom_grid_top_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_4__pin_sc_in_0_(grid_io_bottom_3__1__undriven_top_width_0_height_0_subtile_4__pin_sc_in_0_),
		.top_width_0_height_0_subtile_4__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_4__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_4__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_4__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_4__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_4__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_5__pin_f2a_i_0_(cbx_2__1__1_bottom_grid_top_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_5__pin_sc_in_0_(grid_io_bottom_3__1__undriven_top_width_0_height_0_subtile_5__pin_sc_in_0_),
		.top_width_0_height_0_subtile_5__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_5__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_5__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_5__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_5__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_5__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_6__pin_f2a_i_0_(cbx_2__1__1_bottom_grid_top_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_6__pin_sc_in_0_(grid_io_bottom_3__1__undriven_top_width_0_height_0_subtile_6__pin_sc_in_0_),
		.top_width_0_height_0_subtile_6__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_6__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_6__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_6__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_6__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_6__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_7__pin_f2a_i_0_(cbx_2__1__1_bottom_grid_top_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_7__pin_sc_in_0_(grid_io_bottom_3__1__undriven_top_width_0_height_0_subtile_7__pin_sc_in_0_),
		.top_width_0_height_0_subtile_7__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_7__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_7__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_7__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_7__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_7__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_8__pin_f2a_i_0_(cbx_2__1__1_bottom_grid_top_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_8__pin_sc_in_0_(grid_io_bottom_3__1__undriven_top_width_0_height_0_subtile_8__pin_sc_in_0_),
		.top_width_0_height_0_subtile_8__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_8__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_8__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_8__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_8__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_8__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_9__pin_f2a_i_0_(cbx_2__1__1_bottom_grid_top_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_9__pin_sc_in_0_(grid_io_bottom_3__1__undriven_top_width_0_height_0_subtile_9__pin_sc_in_0_),
		.top_width_0_height_0_subtile_9__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_9__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_9__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_9__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_9__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_9__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_10__pin_f2a_i_0_(cbx_2__1__1_bottom_grid_top_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_10__pin_sc_in_0_(grid_io_bottom_3__1__undriven_top_width_0_height_0_subtile_10__pin_sc_in_0_),
		.top_width_0_height_0_subtile_10__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_10__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_10__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_10__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_10__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_10__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_11__pin_f2a_i_0_(cbx_2__1__1_bottom_grid_top_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_11__pin_sc_in_0_(grid_io_bottom_3__1__undriven_top_width_0_height_0_subtile_11__pin_sc_in_0_),
		.top_width_0_height_0_subtile_11__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_11__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_11__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_11__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_11__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_11__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_12__pin_f2a_i_0_(cbx_2__1__1_bottom_grid_top_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_12__pin_sc_in_0_(grid_io_bottom_3__1__undriven_top_width_0_height_0_subtile_12__pin_sc_in_0_),
		.top_width_0_height_0_subtile_12__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_12__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_12__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_12__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_12__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_12__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_13__pin_f2a_i_0_(cbx_2__1__1_bottom_grid_top_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_13__pin_sc_in_0_(grid_io_bottom_3__1__undriven_top_width_0_height_0_subtile_13__pin_sc_in_0_),
		.top_width_0_height_0_subtile_13__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_13__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_13__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_13__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_13__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_13__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_14__pin_f2a_i_0_(cbx_2__1__1_bottom_grid_top_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_14__pin_sc_in_0_(grid_io_bottom_3__1__undriven_top_width_0_height_0_subtile_14__pin_sc_in_0_),
		.top_width_0_height_0_subtile_14__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_14__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_14__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_14__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_14__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_14__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_15__pin_f2a_i_0_(cbx_2__1__1_bottom_grid_top_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_15__pin_sc_in_0_(grid_io_bottom_3__1__undriven_top_width_0_height_0_subtile_15__pin_sc_in_0_),
		.top_width_0_height_0_subtile_15__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_15__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_15__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_15__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_15__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_15__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_16__pin_f2a_i_0_(cbx_2__1__1_bottom_grid_top_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_16__pin_sc_in_0_(grid_io_bottom_3__1__undriven_top_width_0_height_0_subtile_16__pin_sc_in_0_),
		.top_width_0_height_0_subtile_16__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_16__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_16__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_16__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_16__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_16__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_17__pin_f2a_i_0_(cbx_2__1__1_bottom_grid_top_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_17__pin_sc_in_0_(grid_io_bottom_3__1__undriven_top_width_0_height_0_subtile_17__pin_sc_in_0_),
		.top_width_0_height_0_subtile_17__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_17__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_17__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_17__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_17__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_17__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_18__pin_f2a_i_0_(cbx_2__1__1_bottom_grid_top_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_18__pin_sc_in_0_(grid_io_bottom_3__1__undriven_top_width_0_height_0_subtile_18__pin_sc_in_0_),
		.top_width_0_height_0_subtile_18__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_18__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_18__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_18__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_18__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_18__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_19__pin_f2a_i_0_(cbx_2__1__1_bottom_grid_top_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_19__pin_sc_in_0_(grid_io_bottom_3__1__undriven_top_width_0_height_0_subtile_19__pin_sc_in_0_),
		.top_width_0_height_0_subtile_19__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_19__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_19__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_19__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_19__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_19__pin_clk_3_(clk[3]),
		.ccff_head(sb_2__0__1_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_0__pin_sc_out_0_(grid_io_bottom_3__1__undriven_top_width_0_height_0_subtile_0__pin_sc_out_0_),
		.top_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_1__pin_sc_out_0_(grid_io_bottom_3__1__undriven_top_width_0_height_0_subtile_1__pin_sc_out_0_),
		.top_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_2__pin_sc_out_0_(grid_io_bottom_3__1__undriven_top_width_0_height_0_subtile_2__pin_sc_out_0_),
		.top_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_3__pin_sc_out_0_(grid_io_bottom_3__1__undriven_top_width_0_height_0_subtile_3__pin_sc_out_0_),
		.top_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_4__pin_sc_out_0_(grid_io_bottom_3__1__undriven_top_width_0_height_0_subtile_4__pin_sc_out_0_),
		.top_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_5__pin_sc_out_0_(grid_io_bottom_3__1__undriven_top_width_0_height_0_subtile_5__pin_sc_out_0_),
		.top_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_6__pin_sc_out_0_(grid_io_bottom_3__1__undriven_top_width_0_height_0_subtile_6__pin_sc_out_0_),
		.top_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_7__pin_sc_out_0_(grid_io_bottom_3__1__undriven_top_width_0_height_0_subtile_7__pin_sc_out_0_),
		.top_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_8__pin_sc_out_0_(grid_io_bottom_3__1__undriven_top_width_0_height_0_subtile_8__pin_sc_out_0_),
		.top_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_9__pin_sc_out_0_(grid_io_bottom_3__1__undriven_top_width_0_height_0_subtile_9__pin_sc_out_0_),
		.top_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_10__pin_sc_out_0_(grid_io_bottom_3__1__undriven_top_width_0_height_0_subtile_10__pin_sc_out_0_),
		.top_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_11__pin_sc_out_0_(grid_io_bottom_3__1__undriven_top_width_0_height_0_subtile_11__pin_sc_out_0_),
		.top_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_12__pin_sc_out_0_(grid_io_bottom_3__1__undriven_top_width_0_height_0_subtile_12__pin_sc_out_0_),
		.top_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_13__pin_sc_out_0_(grid_io_bottom_3__1__undriven_top_width_0_height_0_subtile_13__pin_sc_out_0_),
		.top_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_14__pin_sc_out_0_(grid_io_bottom_3__1__undriven_top_width_0_height_0_subtile_14__pin_sc_out_0_),
		.top_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_15__pin_sc_out_0_(grid_io_bottom_3__1__undriven_top_width_0_height_0_subtile_15__pin_sc_out_0_),
		.top_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_16__pin_sc_out_0_(grid_io_bottom_3__1__undriven_top_width_0_height_0_subtile_16__pin_sc_out_0_),
		.top_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_17__pin_sc_out_0_(grid_io_bottom_3__1__undriven_top_width_0_height_0_subtile_17__pin_sc_out_0_),
		.top_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_18__pin_sc_out_0_(grid_io_bottom_3__1__undriven_top_width_0_height_0_subtile_18__pin_sc_out_0_),
		.top_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_19__pin_sc_out_0_(grid_io_bottom_3__1__undriven_top_width_0_height_0_subtile_19__pin_sc_out_0_),
		.ccff_tail(grid_io_bottom_1_ccff_tail));

	grid_io_bottom grid_io_bottom_4__1_ (
		.test_en(test_en),
		.scan_mode(scan_mode),
		.scan_clk(scan_clk),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.CFG_DONE(CFG_DONE),
		.gfpga_pad_QL_PREIO_A2F(gfpga_pad_QL_PREIO_A2F[580:599]),
		.gfpga_pad_QL_PREIO_F2A(gfpga_pad_QL_PREIO_F2A[580:599]),
		.gfpga_pad_QL_PREIO_F2A_DEF0(gfpga_pad_QL_PREIO_F2A_DEF0[580:599]),
		.gfpga_pad_QL_PREIO_F2A_DEF1(gfpga_pad_QL_PREIO_F2A_DEF1[580:599]),
		.gfpga_pad_QL_PREIO_F2A_CLK(gfpga_pad_QL_PREIO_F2A_CLK[580:599]),
		.top_width_0_height_0_subtile_0__pin_f2a_i_0_(cbx_4__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_io_bottom_4__1__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
		.top_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_1__pin_f2a_i_0_(cbx_4__1__0_bottom_grid_top_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_1__pin_sc_in_0_(grid_io_bottom_4__1__undriven_top_width_0_height_0_subtile_1__pin_sc_in_0_),
		.top_width_0_height_0_subtile_1__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_1__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_1__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_1__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_1__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_1__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_2__pin_f2a_i_0_(cbx_4__1__0_bottom_grid_top_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_2__pin_sc_in_0_(grid_io_bottom_4__1__undriven_top_width_0_height_0_subtile_2__pin_sc_in_0_),
		.top_width_0_height_0_subtile_2__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_2__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_2__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_2__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_2__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_2__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_3__pin_f2a_i_0_(cbx_4__1__0_bottom_grid_top_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_3__pin_sc_in_0_(grid_io_bottom_4__1__undriven_top_width_0_height_0_subtile_3__pin_sc_in_0_),
		.top_width_0_height_0_subtile_3__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_3__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_3__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_3__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_3__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_3__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_4__pin_f2a_i_0_(cbx_4__1__0_bottom_grid_top_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_4__pin_sc_in_0_(grid_io_bottom_4__1__undriven_top_width_0_height_0_subtile_4__pin_sc_in_0_),
		.top_width_0_height_0_subtile_4__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_4__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_4__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_4__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_4__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_4__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_5__pin_f2a_i_0_(cbx_4__1__0_bottom_grid_top_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_5__pin_sc_in_0_(grid_io_bottom_4__1__undriven_top_width_0_height_0_subtile_5__pin_sc_in_0_),
		.top_width_0_height_0_subtile_5__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_5__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_5__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_5__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_5__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_5__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_6__pin_f2a_i_0_(cbx_4__1__0_bottom_grid_top_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_6__pin_sc_in_0_(grid_io_bottom_4__1__undriven_top_width_0_height_0_subtile_6__pin_sc_in_0_),
		.top_width_0_height_0_subtile_6__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_6__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_6__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_6__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_6__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_6__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_7__pin_f2a_i_0_(cbx_4__1__0_bottom_grid_top_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_7__pin_sc_in_0_(grid_io_bottom_4__1__undriven_top_width_0_height_0_subtile_7__pin_sc_in_0_),
		.top_width_0_height_0_subtile_7__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_7__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_7__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_7__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_7__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_7__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_8__pin_f2a_i_0_(cbx_4__1__0_bottom_grid_top_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_8__pin_sc_in_0_(grid_io_bottom_4__1__undriven_top_width_0_height_0_subtile_8__pin_sc_in_0_),
		.top_width_0_height_0_subtile_8__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_8__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_8__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_8__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_8__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_8__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_9__pin_f2a_i_0_(cbx_4__1__0_bottom_grid_top_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_9__pin_sc_in_0_(grid_io_bottom_4__1__undriven_top_width_0_height_0_subtile_9__pin_sc_in_0_),
		.top_width_0_height_0_subtile_9__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_9__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_9__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_9__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_9__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_9__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_10__pin_f2a_i_0_(cbx_4__1__0_bottom_grid_top_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_10__pin_sc_in_0_(grid_io_bottom_4__1__undriven_top_width_0_height_0_subtile_10__pin_sc_in_0_),
		.top_width_0_height_0_subtile_10__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_10__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_10__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_10__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_10__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_10__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_11__pin_f2a_i_0_(cbx_4__1__0_bottom_grid_top_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_11__pin_sc_in_0_(grid_io_bottom_4__1__undriven_top_width_0_height_0_subtile_11__pin_sc_in_0_),
		.top_width_0_height_0_subtile_11__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_11__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_11__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_11__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_11__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_11__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_12__pin_f2a_i_0_(cbx_4__1__0_bottom_grid_top_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_12__pin_sc_in_0_(grid_io_bottom_4__1__undriven_top_width_0_height_0_subtile_12__pin_sc_in_0_),
		.top_width_0_height_0_subtile_12__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_12__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_12__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_12__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_12__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_12__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_13__pin_f2a_i_0_(cbx_4__1__0_bottom_grid_top_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_13__pin_sc_in_0_(grid_io_bottom_4__1__undriven_top_width_0_height_0_subtile_13__pin_sc_in_0_),
		.top_width_0_height_0_subtile_13__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_13__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_13__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_13__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_13__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_13__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_14__pin_f2a_i_0_(cbx_4__1__0_bottom_grid_top_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_14__pin_sc_in_0_(grid_io_bottom_4__1__undriven_top_width_0_height_0_subtile_14__pin_sc_in_0_),
		.top_width_0_height_0_subtile_14__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_14__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_14__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_14__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_14__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_14__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_15__pin_f2a_i_0_(cbx_4__1__0_bottom_grid_top_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_15__pin_sc_in_0_(grid_io_bottom_4__1__undriven_top_width_0_height_0_subtile_15__pin_sc_in_0_),
		.top_width_0_height_0_subtile_15__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_15__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_15__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_15__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_15__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_15__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_16__pin_f2a_i_0_(cbx_4__1__0_bottom_grid_top_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_16__pin_sc_in_0_(grid_io_bottom_4__1__undriven_top_width_0_height_0_subtile_16__pin_sc_in_0_),
		.top_width_0_height_0_subtile_16__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_16__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_16__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_16__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_16__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_16__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_17__pin_f2a_i_0_(cbx_4__1__0_bottom_grid_top_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_17__pin_sc_in_0_(grid_io_bottom_4__1__undriven_top_width_0_height_0_subtile_17__pin_sc_in_0_),
		.top_width_0_height_0_subtile_17__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_17__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_17__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_17__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_17__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_17__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_18__pin_f2a_i_0_(cbx_4__1__0_bottom_grid_top_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_18__pin_sc_in_0_(grid_io_bottom_4__1__undriven_top_width_0_height_0_subtile_18__pin_sc_in_0_),
		.top_width_0_height_0_subtile_18__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_18__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_18__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_18__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_18__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_18__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_19__pin_f2a_i_0_(cbx_4__1__0_bottom_grid_top_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_19__pin_sc_in_0_(grid_io_bottom_4__1__undriven_top_width_0_height_0_subtile_19__pin_sc_in_0_),
		.top_width_0_height_0_subtile_19__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_19__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_19__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_19__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_19__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_19__pin_clk_3_(clk[3]),
		.ccff_head(sb_2__0__2_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_0__pin_sc_out_0_(grid_io_bottom_4__1__undriven_top_width_0_height_0_subtile_0__pin_sc_out_0_),
		.top_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_1__pin_sc_out_0_(grid_io_bottom_4__1__undriven_top_width_0_height_0_subtile_1__pin_sc_out_0_),
		.top_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_2__pin_sc_out_0_(grid_io_bottom_4__1__undriven_top_width_0_height_0_subtile_2__pin_sc_out_0_),
		.top_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_3__pin_sc_out_0_(grid_io_bottom_4__1__undriven_top_width_0_height_0_subtile_3__pin_sc_out_0_),
		.top_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_4__pin_sc_out_0_(grid_io_bottom_4__1__undriven_top_width_0_height_0_subtile_4__pin_sc_out_0_),
		.top_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_5__pin_sc_out_0_(grid_io_bottom_4__1__undriven_top_width_0_height_0_subtile_5__pin_sc_out_0_),
		.top_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_6__pin_sc_out_0_(grid_io_bottom_4__1__undriven_top_width_0_height_0_subtile_6__pin_sc_out_0_),
		.top_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_7__pin_sc_out_0_(grid_io_bottom_4__1__undriven_top_width_0_height_0_subtile_7__pin_sc_out_0_),
		.top_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_8__pin_sc_out_0_(grid_io_bottom_4__1__undriven_top_width_0_height_0_subtile_8__pin_sc_out_0_),
		.top_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_9__pin_sc_out_0_(grid_io_bottom_4__1__undriven_top_width_0_height_0_subtile_9__pin_sc_out_0_),
		.top_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_10__pin_sc_out_0_(grid_io_bottom_4__1__undriven_top_width_0_height_0_subtile_10__pin_sc_out_0_),
		.top_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_11__pin_sc_out_0_(grid_io_bottom_4__1__undriven_top_width_0_height_0_subtile_11__pin_sc_out_0_),
		.top_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_12__pin_sc_out_0_(grid_io_bottom_4__1__undriven_top_width_0_height_0_subtile_12__pin_sc_out_0_),
		.top_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_13__pin_sc_out_0_(grid_io_bottom_4__1__undriven_top_width_0_height_0_subtile_13__pin_sc_out_0_),
		.top_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_14__pin_sc_out_0_(grid_io_bottom_4__1__undriven_top_width_0_height_0_subtile_14__pin_sc_out_0_),
		.top_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_15__pin_sc_out_0_(grid_io_bottom_4__1__undriven_top_width_0_height_0_subtile_15__pin_sc_out_0_),
		.top_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_16__pin_sc_out_0_(grid_io_bottom_4__1__undriven_top_width_0_height_0_subtile_16__pin_sc_out_0_),
		.top_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_17__pin_sc_out_0_(grid_io_bottom_4__1__undriven_top_width_0_height_0_subtile_17__pin_sc_out_0_),
		.top_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_18__pin_sc_out_0_(grid_io_bottom_4__1__undriven_top_width_0_height_0_subtile_18__pin_sc_out_0_),
		.top_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_19__pin_sc_out_0_(grid_io_bottom_4__1__undriven_top_width_0_height_0_subtile_19__pin_sc_out_0_),
		.ccff_tail(grid_io_bottom_2_ccff_tail));

	grid_io_bottom grid_io_bottom_5__1_ (
		.test_en(test_en),
		.scan_mode(scan_mode),
		.scan_clk(scan_clk),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.CFG_DONE(CFG_DONE),
		.gfpga_pad_QL_PREIO_A2F(gfpga_pad_QL_PREIO_A2F[560:579]),
		.gfpga_pad_QL_PREIO_F2A(gfpga_pad_QL_PREIO_F2A[560:579]),
		.gfpga_pad_QL_PREIO_F2A_DEF0(gfpga_pad_QL_PREIO_F2A_DEF0[560:579]),
		.gfpga_pad_QL_PREIO_F2A_DEF1(gfpga_pad_QL_PREIO_F2A_DEF1[560:579]),
		.gfpga_pad_QL_PREIO_F2A_CLK(gfpga_pad_QL_PREIO_F2A_CLK[560:579]),
		.top_width_0_height_0_subtile_0__pin_f2a_i_0_(cbx_2__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_io_bottom_5__1__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
		.top_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_1__pin_f2a_i_0_(cbx_2__1__2_bottom_grid_top_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_1__pin_sc_in_0_(grid_io_bottom_5__1__undriven_top_width_0_height_0_subtile_1__pin_sc_in_0_),
		.top_width_0_height_0_subtile_1__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_1__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_1__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_1__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_1__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_1__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_2__pin_f2a_i_0_(cbx_2__1__2_bottom_grid_top_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_2__pin_sc_in_0_(grid_io_bottom_5__1__undriven_top_width_0_height_0_subtile_2__pin_sc_in_0_),
		.top_width_0_height_0_subtile_2__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_2__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_2__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_2__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_2__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_2__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_3__pin_f2a_i_0_(cbx_2__1__2_bottom_grid_top_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_3__pin_sc_in_0_(grid_io_bottom_5__1__undriven_top_width_0_height_0_subtile_3__pin_sc_in_0_),
		.top_width_0_height_0_subtile_3__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_3__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_3__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_3__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_3__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_3__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_4__pin_f2a_i_0_(cbx_2__1__2_bottom_grid_top_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_4__pin_sc_in_0_(grid_io_bottom_5__1__undriven_top_width_0_height_0_subtile_4__pin_sc_in_0_),
		.top_width_0_height_0_subtile_4__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_4__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_4__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_4__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_4__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_4__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_5__pin_f2a_i_0_(cbx_2__1__2_bottom_grid_top_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_5__pin_sc_in_0_(grid_io_bottom_5__1__undriven_top_width_0_height_0_subtile_5__pin_sc_in_0_),
		.top_width_0_height_0_subtile_5__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_5__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_5__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_5__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_5__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_5__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_6__pin_f2a_i_0_(cbx_2__1__2_bottom_grid_top_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_6__pin_sc_in_0_(grid_io_bottom_5__1__undriven_top_width_0_height_0_subtile_6__pin_sc_in_0_),
		.top_width_0_height_0_subtile_6__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_6__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_6__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_6__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_6__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_6__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_7__pin_f2a_i_0_(cbx_2__1__2_bottom_grid_top_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_7__pin_sc_in_0_(grid_io_bottom_5__1__undriven_top_width_0_height_0_subtile_7__pin_sc_in_0_),
		.top_width_0_height_0_subtile_7__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_7__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_7__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_7__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_7__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_7__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_8__pin_f2a_i_0_(cbx_2__1__2_bottom_grid_top_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_8__pin_sc_in_0_(grid_io_bottom_5__1__undriven_top_width_0_height_0_subtile_8__pin_sc_in_0_),
		.top_width_0_height_0_subtile_8__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_8__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_8__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_8__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_8__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_8__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_9__pin_f2a_i_0_(cbx_2__1__2_bottom_grid_top_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_9__pin_sc_in_0_(grid_io_bottom_5__1__undriven_top_width_0_height_0_subtile_9__pin_sc_in_0_),
		.top_width_0_height_0_subtile_9__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_9__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_9__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_9__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_9__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_9__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_10__pin_f2a_i_0_(cbx_2__1__2_bottom_grid_top_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_10__pin_sc_in_0_(grid_io_bottom_5__1__undriven_top_width_0_height_0_subtile_10__pin_sc_in_0_),
		.top_width_0_height_0_subtile_10__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_10__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_10__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_10__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_10__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_10__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_11__pin_f2a_i_0_(cbx_2__1__2_bottom_grid_top_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_11__pin_sc_in_0_(grid_io_bottom_5__1__undriven_top_width_0_height_0_subtile_11__pin_sc_in_0_),
		.top_width_0_height_0_subtile_11__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_11__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_11__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_11__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_11__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_11__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_12__pin_f2a_i_0_(cbx_2__1__2_bottom_grid_top_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_12__pin_sc_in_0_(grid_io_bottom_5__1__undriven_top_width_0_height_0_subtile_12__pin_sc_in_0_),
		.top_width_0_height_0_subtile_12__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_12__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_12__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_12__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_12__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_12__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_13__pin_f2a_i_0_(cbx_2__1__2_bottom_grid_top_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_13__pin_sc_in_0_(grid_io_bottom_5__1__undriven_top_width_0_height_0_subtile_13__pin_sc_in_0_),
		.top_width_0_height_0_subtile_13__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_13__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_13__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_13__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_13__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_13__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_14__pin_f2a_i_0_(cbx_2__1__2_bottom_grid_top_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_14__pin_sc_in_0_(grid_io_bottom_5__1__undriven_top_width_0_height_0_subtile_14__pin_sc_in_0_),
		.top_width_0_height_0_subtile_14__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_14__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_14__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_14__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_14__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_14__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_15__pin_f2a_i_0_(cbx_2__1__2_bottom_grid_top_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_15__pin_sc_in_0_(grid_io_bottom_5__1__undriven_top_width_0_height_0_subtile_15__pin_sc_in_0_),
		.top_width_0_height_0_subtile_15__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_15__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_15__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_15__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_15__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_15__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_16__pin_f2a_i_0_(cbx_2__1__2_bottom_grid_top_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_16__pin_sc_in_0_(grid_io_bottom_5__1__undriven_top_width_0_height_0_subtile_16__pin_sc_in_0_),
		.top_width_0_height_0_subtile_16__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_16__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_16__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_16__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_16__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_16__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_17__pin_f2a_i_0_(cbx_2__1__2_bottom_grid_top_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_17__pin_sc_in_0_(grid_io_bottom_5__1__undriven_top_width_0_height_0_subtile_17__pin_sc_in_0_),
		.top_width_0_height_0_subtile_17__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_17__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_17__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_17__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_17__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_17__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_18__pin_f2a_i_0_(cbx_2__1__2_bottom_grid_top_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_18__pin_sc_in_0_(grid_io_bottom_5__1__undriven_top_width_0_height_0_subtile_18__pin_sc_in_0_),
		.top_width_0_height_0_subtile_18__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_18__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_18__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_18__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_18__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_18__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_19__pin_f2a_i_0_(cbx_2__1__2_bottom_grid_top_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_19__pin_sc_in_0_(grid_io_bottom_5__1__undriven_top_width_0_height_0_subtile_19__pin_sc_in_0_),
		.top_width_0_height_0_subtile_19__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_19__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_19__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_19__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_19__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_19__pin_clk_3_(clk[3]),
		.ccff_head(sb_2__0__3_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_0__pin_sc_out_0_(grid_io_bottom_5__1__undriven_top_width_0_height_0_subtile_0__pin_sc_out_0_),
		.top_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_1__pin_sc_out_0_(grid_io_bottom_5__1__undriven_top_width_0_height_0_subtile_1__pin_sc_out_0_),
		.top_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_2__pin_sc_out_0_(grid_io_bottom_5__1__undriven_top_width_0_height_0_subtile_2__pin_sc_out_0_),
		.top_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_3__pin_sc_out_0_(grid_io_bottom_5__1__undriven_top_width_0_height_0_subtile_3__pin_sc_out_0_),
		.top_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_4__pin_sc_out_0_(grid_io_bottom_5__1__undriven_top_width_0_height_0_subtile_4__pin_sc_out_0_),
		.top_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_5__pin_sc_out_0_(grid_io_bottom_5__1__undriven_top_width_0_height_0_subtile_5__pin_sc_out_0_),
		.top_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_6__pin_sc_out_0_(grid_io_bottom_5__1__undriven_top_width_0_height_0_subtile_6__pin_sc_out_0_),
		.top_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_7__pin_sc_out_0_(grid_io_bottom_5__1__undriven_top_width_0_height_0_subtile_7__pin_sc_out_0_),
		.top_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_8__pin_sc_out_0_(grid_io_bottom_5__1__undriven_top_width_0_height_0_subtile_8__pin_sc_out_0_),
		.top_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_9__pin_sc_out_0_(grid_io_bottom_5__1__undriven_top_width_0_height_0_subtile_9__pin_sc_out_0_),
		.top_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_10__pin_sc_out_0_(grid_io_bottom_5__1__undriven_top_width_0_height_0_subtile_10__pin_sc_out_0_),
		.top_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_11__pin_sc_out_0_(grid_io_bottom_5__1__undriven_top_width_0_height_0_subtile_11__pin_sc_out_0_),
		.top_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_12__pin_sc_out_0_(grid_io_bottom_5__1__undriven_top_width_0_height_0_subtile_12__pin_sc_out_0_),
		.top_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_13__pin_sc_out_0_(grid_io_bottom_5__1__undriven_top_width_0_height_0_subtile_13__pin_sc_out_0_),
		.top_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_14__pin_sc_out_0_(grid_io_bottom_5__1__undriven_top_width_0_height_0_subtile_14__pin_sc_out_0_),
		.top_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_15__pin_sc_out_0_(grid_io_bottom_5__1__undriven_top_width_0_height_0_subtile_15__pin_sc_out_0_),
		.top_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_16__pin_sc_out_0_(grid_io_bottom_5__1__undriven_top_width_0_height_0_subtile_16__pin_sc_out_0_),
		.top_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_17__pin_sc_out_0_(grid_io_bottom_5__1__undriven_top_width_0_height_0_subtile_17__pin_sc_out_0_),
		.top_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_18__pin_sc_out_0_(grid_io_bottom_5__1__undriven_top_width_0_height_0_subtile_18__pin_sc_out_0_),
		.top_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_19__pin_sc_out_0_(grid_io_bottom_5__1__undriven_top_width_0_height_0_subtile_19__pin_sc_out_0_),
		.ccff_tail(ccff_tail[0]));

	grid_io_bottom grid_io_bottom_6__1_ (
		.test_en(test_en),
		.scan_mode(scan_mode),
		.scan_clk(scan_clk),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.CFG_DONE(CFG_DONE),
		.gfpga_pad_QL_PREIO_A2F(gfpga_pad_QL_PREIO_A2F[540:559]),
		.gfpga_pad_QL_PREIO_F2A(gfpga_pad_QL_PREIO_F2A[540:559]),
		.gfpga_pad_QL_PREIO_F2A_DEF0(gfpga_pad_QL_PREIO_F2A_DEF0[540:559]),
		.gfpga_pad_QL_PREIO_F2A_DEF1(gfpga_pad_QL_PREIO_F2A_DEF1[540:559]),
		.gfpga_pad_QL_PREIO_F2A_CLK(gfpga_pad_QL_PREIO_F2A_CLK[540:559]),
		.top_width_0_height_0_subtile_0__pin_f2a_i_0_(cbx_2__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_io_bottom_6__1__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
		.top_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_1__pin_f2a_i_0_(cbx_2__1__3_bottom_grid_top_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_1__pin_sc_in_0_(grid_io_bottom_6__1__undriven_top_width_0_height_0_subtile_1__pin_sc_in_0_),
		.top_width_0_height_0_subtile_1__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_1__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_1__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_1__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_1__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_1__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_2__pin_f2a_i_0_(cbx_2__1__3_bottom_grid_top_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_2__pin_sc_in_0_(grid_io_bottom_6__1__undriven_top_width_0_height_0_subtile_2__pin_sc_in_0_),
		.top_width_0_height_0_subtile_2__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_2__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_2__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_2__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_2__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_2__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_3__pin_f2a_i_0_(cbx_2__1__3_bottom_grid_top_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_3__pin_sc_in_0_(grid_io_bottom_6__1__undriven_top_width_0_height_0_subtile_3__pin_sc_in_0_),
		.top_width_0_height_0_subtile_3__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_3__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_3__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_3__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_3__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_3__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_4__pin_f2a_i_0_(cbx_2__1__3_bottom_grid_top_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_4__pin_sc_in_0_(grid_io_bottom_6__1__undriven_top_width_0_height_0_subtile_4__pin_sc_in_0_),
		.top_width_0_height_0_subtile_4__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_4__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_4__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_4__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_4__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_4__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_5__pin_f2a_i_0_(cbx_2__1__3_bottom_grid_top_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_5__pin_sc_in_0_(grid_io_bottom_6__1__undriven_top_width_0_height_0_subtile_5__pin_sc_in_0_),
		.top_width_0_height_0_subtile_5__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_5__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_5__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_5__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_5__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_5__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_6__pin_f2a_i_0_(cbx_2__1__3_bottom_grid_top_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_6__pin_sc_in_0_(grid_io_bottom_6__1__undriven_top_width_0_height_0_subtile_6__pin_sc_in_0_),
		.top_width_0_height_0_subtile_6__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_6__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_6__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_6__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_6__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_6__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_7__pin_f2a_i_0_(cbx_2__1__3_bottom_grid_top_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_7__pin_sc_in_0_(grid_io_bottom_6__1__undriven_top_width_0_height_0_subtile_7__pin_sc_in_0_),
		.top_width_0_height_0_subtile_7__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_7__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_7__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_7__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_7__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_7__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_8__pin_f2a_i_0_(cbx_2__1__3_bottom_grid_top_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_8__pin_sc_in_0_(grid_io_bottom_6__1__undriven_top_width_0_height_0_subtile_8__pin_sc_in_0_),
		.top_width_0_height_0_subtile_8__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_8__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_8__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_8__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_8__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_8__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_9__pin_f2a_i_0_(cbx_2__1__3_bottom_grid_top_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_9__pin_sc_in_0_(grid_io_bottom_6__1__undriven_top_width_0_height_0_subtile_9__pin_sc_in_0_),
		.top_width_0_height_0_subtile_9__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_9__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_9__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_9__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_9__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_9__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_10__pin_f2a_i_0_(cbx_2__1__3_bottom_grid_top_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_10__pin_sc_in_0_(grid_io_bottom_6__1__undriven_top_width_0_height_0_subtile_10__pin_sc_in_0_),
		.top_width_0_height_0_subtile_10__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_10__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_10__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_10__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_10__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_10__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_11__pin_f2a_i_0_(cbx_2__1__3_bottom_grid_top_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_11__pin_sc_in_0_(grid_io_bottom_6__1__undriven_top_width_0_height_0_subtile_11__pin_sc_in_0_),
		.top_width_0_height_0_subtile_11__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_11__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_11__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_11__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_11__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_11__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_12__pin_f2a_i_0_(cbx_2__1__3_bottom_grid_top_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_12__pin_sc_in_0_(grid_io_bottom_6__1__undriven_top_width_0_height_0_subtile_12__pin_sc_in_0_),
		.top_width_0_height_0_subtile_12__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_12__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_12__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_12__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_12__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_12__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_13__pin_f2a_i_0_(cbx_2__1__3_bottom_grid_top_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_13__pin_sc_in_0_(grid_io_bottom_6__1__undriven_top_width_0_height_0_subtile_13__pin_sc_in_0_),
		.top_width_0_height_0_subtile_13__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_13__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_13__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_13__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_13__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_13__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_14__pin_f2a_i_0_(cbx_2__1__3_bottom_grid_top_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_14__pin_sc_in_0_(grid_io_bottom_6__1__undriven_top_width_0_height_0_subtile_14__pin_sc_in_0_),
		.top_width_0_height_0_subtile_14__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_14__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_14__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_14__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_14__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_14__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_15__pin_f2a_i_0_(cbx_2__1__3_bottom_grid_top_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_15__pin_sc_in_0_(grid_io_bottom_6__1__undriven_top_width_0_height_0_subtile_15__pin_sc_in_0_),
		.top_width_0_height_0_subtile_15__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_15__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_15__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_15__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_15__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_15__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_16__pin_f2a_i_0_(cbx_2__1__3_bottom_grid_top_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_16__pin_sc_in_0_(grid_io_bottom_6__1__undriven_top_width_0_height_0_subtile_16__pin_sc_in_0_),
		.top_width_0_height_0_subtile_16__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_16__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_16__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_16__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_16__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_16__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_17__pin_f2a_i_0_(cbx_2__1__3_bottom_grid_top_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_17__pin_sc_in_0_(grid_io_bottom_6__1__undriven_top_width_0_height_0_subtile_17__pin_sc_in_0_),
		.top_width_0_height_0_subtile_17__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_17__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_17__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_17__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_17__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_17__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_18__pin_f2a_i_0_(cbx_2__1__3_bottom_grid_top_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_18__pin_sc_in_0_(grid_io_bottom_6__1__undriven_top_width_0_height_0_subtile_18__pin_sc_in_0_),
		.top_width_0_height_0_subtile_18__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_18__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_18__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_18__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_18__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_18__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_19__pin_f2a_i_0_(cbx_2__1__3_bottom_grid_top_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_19__pin_sc_in_0_(grid_io_bottom_6__1__undriven_top_width_0_height_0_subtile_19__pin_sc_in_0_),
		.top_width_0_height_0_subtile_19__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_19__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_19__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_19__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_19__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_19__pin_clk_3_(clk[3]),
		.ccff_head(sb_2__0__4_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_0__pin_sc_out_0_(grid_io_bottom_6__1__undriven_top_width_0_height_0_subtile_0__pin_sc_out_0_),
		.top_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_1__pin_sc_out_0_(grid_io_bottom_6__1__undriven_top_width_0_height_0_subtile_1__pin_sc_out_0_),
		.top_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_2__pin_sc_out_0_(grid_io_bottom_6__1__undriven_top_width_0_height_0_subtile_2__pin_sc_out_0_),
		.top_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_3__pin_sc_out_0_(grid_io_bottom_6__1__undriven_top_width_0_height_0_subtile_3__pin_sc_out_0_),
		.top_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_4__pin_sc_out_0_(grid_io_bottom_6__1__undriven_top_width_0_height_0_subtile_4__pin_sc_out_0_),
		.top_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_5__pin_sc_out_0_(grid_io_bottom_6__1__undriven_top_width_0_height_0_subtile_5__pin_sc_out_0_),
		.top_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_6__pin_sc_out_0_(grid_io_bottom_6__1__undriven_top_width_0_height_0_subtile_6__pin_sc_out_0_),
		.top_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_7__pin_sc_out_0_(grid_io_bottom_6__1__undriven_top_width_0_height_0_subtile_7__pin_sc_out_0_),
		.top_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_8__pin_sc_out_0_(grid_io_bottom_6__1__undriven_top_width_0_height_0_subtile_8__pin_sc_out_0_),
		.top_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_9__pin_sc_out_0_(grid_io_bottom_6__1__undriven_top_width_0_height_0_subtile_9__pin_sc_out_0_),
		.top_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_10__pin_sc_out_0_(grid_io_bottom_6__1__undriven_top_width_0_height_0_subtile_10__pin_sc_out_0_),
		.top_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_11__pin_sc_out_0_(grid_io_bottom_6__1__undriven_top_width_0_height_0_subtile_11__pin_sc_out_0_),
		.top_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_12__pin_sc_out_0_(grid_io_bottom_6__1__undriven_top_width_0_height_0_subtile_12__pin_sc_out_0_),
		.top_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_13__pin_sc_out_0_(grid_io_bottom_6__1__undriven_top_width_0_height_0_subtile_13__pin_sc_out_0_),
		.top_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_14__pin_sc_out_0_(grid_io_bottom_6__1__undriven_top_width_0_height_0_subtile_14__pin_sc_out_0_),
		.top_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_15__pin_sc_out_0_(grid_io_bottom_6__1__undriven_top_width_0_height_0_subtile_15__pin_sc_out_0_),
		.top_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_16__pin_sc_out_0_(grid_io_bottom_6__1__undriven_top_width_0_height_0_subtile_16__pin_sc_out_0_),
		.top_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_17__pin_sc_out_0_(grid_io_bottom_6__1__undriven_top_width_0_height_0_subtile_17__pin_sc_out_0_),
		.top_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_18__pin_sc_out_0_(grid_io_bottom_6__1__undriven_top_width_0_height_0_subtile_18__pin_sc_out_0_),
		.top_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_19__pin_sc_out_0_(grid_io_bottom_6__1__undriven_top_width_0_height_0_subtile_19__pin_sc_out_0_),
		.ccff_tail(grid_io_bottom_4_ccff_tail));

	grid_io_bottom grid_io_bottom_7__1_ (
		.test_en(test_en),
		.scan_mode(scan_mode),
		.scan_clk(scan_clk),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.CFG_DONE(CFG_DONE),
		.gfpga_pad_QL_PREIO_A2F(gfpga_pad_QL_PREIO_A2F[520:539]),
		.gfpga_pad_QL_PREIO_F2A(gfpga_pad_QL_PREIO_F2A[520:539]),
		.gfpga_pad_QL_PREIO_F2A_DEF0(gfpga_pad_QL_PREIO_F2A_DEF0[520:539]),
		.gfpga_pad_QL_PREIO_F2A_DEF1(gfpga_pad_QL_PREIO_F2A_DEF1[520:539]),
		.gfpga_pad_QL_PREIO_F2A_CLK(gfpga_pad_QL_PREIO_F2A_CLK[520:539]),
		.top_width_0_height_0_subtile_0__pin_f2a_i_0_(cbx_7__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_io_bottom_7__1__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
		.top_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_1__pin_f2a_i_0_(cbx_7__1__0_bottom_grid_top_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_1__pin_sc_in_0_(grid_io_bottom_7__1__undriven_top_width_0_height_0_subtile_1__pin_sc_in_0_),
		.top_width_0_height_0_subtile_1__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_1__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_1__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_1__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_1__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_1__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_2__pin_f2a_i_0_(cbx_7__1__0_bottom_grid_top_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_2__pin_sc_in_0_(grid_io_bottom_7__1__undriven_top_width_0_height_0_subtile_2__pin_sc_in_0_),
		.top_width_0_height_0_subtile_2__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_2__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_2__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_2__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_2__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_2__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_3__pin_f2a_i_0_(cbx_7__1__0_bottom_grid_top_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_3__pin_sc_in_0_(grid_io_bottom_7__1__undriven_top_width_0_height_0_subtile_3__pin_sc_in_0_),
		.top_width_0_height_0_subtile_3__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_3__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_3__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_3__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_3__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_3__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_4__pin_f2a_i_0_(cbx_7__1__0_bottom_grid_top_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_4__pin_sc_in_0_(grid_io_bottom_7__1__undriven_top_width_0_height_0_subtile_4__pin_sc_in_0_),
		.top_width_0_height_0_subtile_4__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_4__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_4__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_4__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_4__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_4__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_5__pin_f2a_i_0_(cbx_7__1__0_bottom_grid_top_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_5__pin_sc_in_0_(grid_io_bottom_7__1__undriven_top_width_0_height_0_subtile_5__pin_sc_in_0_),
		.top_width_0_height_0_subtile_5__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_5__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_5__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_5__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_5__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_5__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_6__pin_f2a_i_0_(cbx_7__1__0_bottom_grid_top_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_6__pin_sc_in_0_(grid_io_bottom_7__1__undriven_top_width_0_height_0_subtile_6__pin_sc_in_0_),
		.top_width_0_height_0_subtile_6__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_6__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_6__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_6__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_6__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_6__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_7__pin_f2a_i_0_(cbx_7__1__0_bottom_grid_top_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_7__pin_sc_in_0_(grid_io_bottom_7__1__undriven_top_width_0_height_0_subtile_7__pin_sc_in_0_),
		.top_width_0_height_0_subtile_7__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_7__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_7__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_7__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_7__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_7__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_8__pin_f2a_i_0_(cbx_7__1__0_bottom_grid_top_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_8__pin_sc_in_0_(grid_io_bottom_7__1__undriven_top_width_0_height_0_subtile_8__pin_sc_in_0_),
		.top_width_0_height_0_subtile_8__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_8__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_8__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_8__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_8__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_8__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_9__pin_f2a_i_0_(cbx_7__1__0_bottom_grid_top_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_9__pin_sc_in_0_(grid_io_bottom_7__1__undriven_top_width_0_height_0_subtile_9__pin_sc_in_0_),
		.top_width_0_height_0_subtile_9__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_9__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_9__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_9__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_9__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_9__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_10__pin_f2a_i_0_(cbx_7__1__0_bottom_grid_top_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_10__pin_sc_in_0_(grid_io_bottom_7__1__undriven_top_width_0_height_0_subtile_10__pin_sc_in_0_),
		.top_width_0_height_0_subtile_10__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_10__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_10__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_10__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_10__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_10__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_11__pin_f2a_i_0_(cbx_7__1__0_bottom_grid_top_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_11__pin_sc_in_0_(grid_io_bottom_7__1__undriven_top_width_0_height_0_subtile_11__pin_sc_in_0_),
		.top_width_0_height_0_subtile_11__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_11__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_11__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_11__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_11__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_11__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_12__pin_f2a_i_0_(cbx_7__1__0_bottom_grid_top_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_12__pin_sc_in_0_(grid_io_bottom_7__1__undriven_top_width_0_height_0_subtile_12__pin_sc_in_0_),
		.top_width_0_height_0_subtile_12__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_12__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_12__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_12__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_12__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_12__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_13__pin_f2a_i_0_(cbx_7__1__0_bottom_grid_top_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_13__pin_sc_in_0_(grid_io_bottom_7__1__undriven_top_width_0_height_0_subtile_13__pin_sc_in_0_),
		.top_width_0_height_0_subtile_13__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_13__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_13__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_13__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_13__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_13__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_14__pin_f2a_i_0_(cbx_7__1__0_bottom_grid_top_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_14__pin_sc_in_0_(grid_io_bottom_7__1__undriven_top_width_0_height_0_subtile_14__pin_sc_in_0_),
		.top_width_0_height_0_subtile_14__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_14__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_14__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_14__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_14__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_14__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_15__pin_f2a_i_0_(cbx_7__1__0_bottom_grid_top_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_15__pin_sc_in_0_(grid_io_bottom_7__1__undriven_top_width_0_height_0_subtile_15__pin_sc_in_0_),
		.top_width_0_height_0_subtile_15__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_15__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_15__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_15__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_15__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_15__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_16__pin_f2a_i_0_(cbx_7__1__0_bottom_grid_top_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_16__pin_sc_in_0_(grid_io_bottom_7__1__undriven_top_width_0_height_0_subtile_16__pin_sc_in_0_),
		.top_width_0_height_0_subtile_16__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_16__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_16__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_16__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_16__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_16__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_17__pin_f2a_i_0_(cbx_7__1__0_bottom_grid_top_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_17__pin_sc_in_0_(grid_io_bottom_7__1__undriven_top_width_0_height_0_subtile_17__pin_sc_in_0_),
		.top_width_0_height_0_subtile_17__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_17__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_17__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_17__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_17__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_17__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_18__pin_f2a_i_0_(cbx_7__1__0_bottom_grid_top_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_18__pin_sc_in_0_(grid_io_bottom_7__1__undriven_top_width_0_height_0_subtile_18__pin_sc_in_0_),
		.top_width_0_height_0_subtile_18__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_18__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_18__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_18__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_18__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_18__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_19__pin_f2a_i_0_(cbx_7__1__0_bottom_grid_top_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_19__pin_sc_in_0_(grid_io_bottom_7__1__undriven_top_width_0_height_0_subtile_19__pin_sc_in_0_),
		.top_width_0_height_0_subtile_19__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_19__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_19__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_19__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_19__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_19__pin_clk_3_(clk[3]),
		.ccff_head(sb_2__0__5_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_0__pin_sc_out_0_(grid_io_bottom_7__1__undriven_top_width_0_height_0_subtile_0__pin_sc_out_0_),
		.top_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_1__pin_sc_out_0_(grid_io_bottom_7__1__undriven_top_width_0_height_0_subtile_1__pin_sc_out_0_),
		.top_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_2__pin_sc_out_0_(grid_io_bottom_7__1__undriven_top_width_0_height_0_subtile_2__pin_sc_out_0_),
		.top_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_3__pin_sc_out_0_(grid_io_bottom_7__1__undriven_top_width_0_height_0_subtile_3__pin_sc_out_0_),
		.top_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_4__pin_sc_out_0_(grid_io_bottom_7__1__undriven_top_width_0_height_0_subtile_4__pin_sc_out_0_),
		.top_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_5__pin_sc_out_0_(grid_io_bottom_7__1__undriven_top_width_0_height_0_subtile_5__pin_sc_out_0_),
		.top_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_6__pin_sc_out_0_(grid_io_bottom_7__1__undriven_top_width_0_height_0_subtile_6__pin_sc_out_0_),
		.top_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_7__pin_sc_out_0_(grid_io_bottom_7__1__undriven_top_width_0_height_0_subtile_7__pin_sc_out_0_),
		.top_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_8__pin_sc_out_0_(grid_io_bottom_7__1__undriven_top_width_0_height_0_subtile_8__pin_sc_out_0_),
		.top_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_9__pin_sc_out_0_(grid_io_bottom_7__1__undriven_top_width_0_height_0_subtile_9__pin_sc_out_0_),
		.top_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_10__pin_sc_out_0_(grid_io_bottom_7__1__undriven_top_width_0_height_0_subtile_10__pin_sc_out_0_),
		.top_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_11__pin_sc_out_0_(grid_io_bottom_7__1__undriven_top_width_0_height_0_subtile_11__pin_sc_out_0_),
		.top_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_12__pin_sc_out_0_(grid_io_bottom_7__1__undriven_top_width_0_height_0_subtile_12__pin_sc_out_0_),
		.top_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_13__pin_sc_out_0_(grid_io_bottom_7__1__undriven_top_width_0_height_0_subtile_13__pin_sc_out_0_),
		.top_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_14__pin_sc_out_0_(grid_io_bottom_7__1__undriven_top_width_0_height_0_subtile_14__pin_sc_out_0_),
		.top_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_15__pin_sc_out_0_(grid_io_bottom_7__1__undriven_top_width_0_height_0_subtile_15__pin_sc_out_0_),
		.top_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_16__pin_sc_out_0_(grid_io_bottom_7__1__undriven_top_width_0_height_0_subtile_16__pin_sc_out_0_),
		.top_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_17__pin_sc_out_0_(grid_io_bottom_7__1__undriven_top_width_0_height_0_subtile_17__pin_sc_out_0_),
		.top_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_18__pin_sc_out_0_(grid_io_bottom_7__1__undriven_top_width_0_height_0_subtile_18__pin_sc_out_0_),
		.top_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_19__pin_sc_out_0_(grid_io_bottom_7__1__undriven_top_width_0_height_0_subtile_19__pin_sc_out_0_),
		.ccff_tail(grid_io_bottom_5_ccff_tail));

	grid_io_bottom grid_io_bottom_8__1_ (
		.test_en(test_en),
		.scan_mode(scan_mode),
		.scan_clk(scan_clk),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.CFG_DONE(CFG_DONE),
		.gfpga_pad_QL_PREIO_A2F(gfpga_pad_QL_PREIO_A2F[500:519]),
		.gfpga_pad_QL_PREIO_F2A(gfpga_pad_QL_PREIO_F2A[500:519]),
		.gfpga_pad_QL_PREIO_F2A_DEF0(gfpga_pad_QL_PREIO_F2A_DEF0[500:519]),
		.gfpga_pad_QL_PREIO_F2A_DEF1(gfpga_pad_QL_PREIO_F2A_DEF1[500:519]),
		.gfpga_pad_QL_PREIO_F2A_CLK(gfpga_pad_QL_PREIO_F2A_CLK[500:519]),
		.top_width_0_height_0_subtile_0__pin_f2a_i_0_(cbx_2__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_io_bottom_8__1__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
		.top_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_1__pin_f2a_i_0_(cbx_2__1__4_bottom_grid_top_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_1__pin_sc_in_0_(grid_io_bottom_8__1__undriven_top_width_0_height_0_subtile_1__pin_sc_in_0_),
		.top_width_0_height_0_subtile_1__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_1__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_1__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_1__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_1__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_1__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_2__pin_f2a_i_0_(cbx_2__1__4_bottom_grid_top_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_2__pin_sc_in_0_(grid_io_bottom_8__1__undriven_top_width_0_height_0_subtile_2__pin_sc_in_0_),
		.top_width_0_height_0_subtile_2__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_2__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_2__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_2__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_2__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_2__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_3__pin_f2a_i_0_(cbx_2__1__4_bottom_grid_top_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_3__pin_sc_in_0_(grid_io_bottom_8__1__undriven_top_width_0_height_0_subtile_3__pin_sc_in_0_),
		.top_width_0_height_0_subtile_3__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_3__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_3__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_3__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_3__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_3__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_4__pin_f2a_i_0_(cbx_2__1__4_bottom_grid_top_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_4__pin_sc_in_0_(grid_io_bottom_8__1__undriven_top_width_0_height_0_subtile_4__pin_sc_in_0_),
		.top_width_0_height_0_subtile_4__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_4__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_4__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_4__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_4__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_4__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_5__pin_f2a_i_0_(cbx_2__1__4_bottom_grid_top_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_5__pin_sc_in_0_(grid_io_bottom_8__1__undriven_top_width_0_height_0_subtile_5__pin_sc_in_0_),
		.top_width_0_height_0_subtile_5__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_5__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_5__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_5__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_5__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_5__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_6__pin_f2a_i_0_(cbx_2__1__4_bottom_grid_top_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_6__pin_sc_in_0_(grid_io_bottom_8__1__undriven_top_width_0_height_0_subtile_6__pin_sc_in_0_),
		.top_width_0_height_0_subtile_6__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_6__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_6__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_6__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_6__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_6__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_7__pin_f2a_i_0_(cbx_2__1__4_bottom_grid_top_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_7__pin_sc_in_0_(grid_io_bottom_8__1__undriven_top_width_0_height_0_subtile_7__pin_sc_in_0_),
		.top_width_0_height_0_subtile_7__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_7__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_7__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_7__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_7__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_7__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_8__pin_f2a_i_0_(cbx_2__1__4_bottom_grid_top_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_8__pin_sc_in_0_(grid_io_bottom_8__1__undriven_top_width_0_height_0_subtile_8__pin_sc_in_0_),
		.top_width_0_height_0_subtile_8__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_8__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_8__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_8__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_8__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_8__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_9__pin_f2a_i_0_(cbx_2__1__4_bottom_grid_top_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_9__pin_sc_in_0_(grid_io_bottom_8__1__undriven_top_width_0_height_0_subtile_9__pin_sc_in_0_),
		.top_width_0_height_0_subtile_9__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_9__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_9__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_9__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_9__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_9__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_10__pin_f2a_i_0_(cbx_2__1__4_bottom_grid_top_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_10__pin_sc_in_0_(grid_io_bottom_8__1__undriven_top_width_0_height_0_subtile_10__pin_sc_in_0_),
		.top_width_0_height_0_subtile_10__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_10__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_10__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_10__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_10__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_10__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_11__pin_f2a_i_0_(cbx_2__1__4_bottom_grid_top_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_11__pin_sc_in_0_(grid_io_bottom_8__1__undriven_top_width_0_height_0_subtile_11__pin_sc_in_0_),
		.top_width_0_height_0_subtile_11__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_11__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_11__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_11__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_11__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_11__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_12__pin_f2a_i_0_(cbx_2__1__4_bottom_grid_top_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_12__pin_sc_in_0_(grid_io_bottom_8__1__undriven_top_width_0_height_0_subtile_12__pin_sc_in_0_),
		.top_width_0_height_0_subtile_12__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_12__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_12__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_12__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_12__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_12__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_13__pin_f2a_i_0_(cbx_2__1__4_bottom_grid_top_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_13__pin_sc_in_0_(grid_io_bottom_8__1__undriven_top_width_0_height_0_subtile_13__pin_sc_in_0_),
		.top_width_0_height_0_subtile_13__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_13__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_13__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_13__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_13__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_13__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_14__pin_f2a_i_0_(cbx_2__1__4_bottom_grid_top_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_14__pin_sc_in_0_(grid_io_bottom_8__1__undriven_top_width_0_height_0_subtile_14__pin_sc_in_0_),
		.top_width_0_height_0_subtile_14__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_14__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_14__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_14__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_14__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_14__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_15__pin_f2a_i_0_(cbx_2__1__4_bottom_grid_top_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_15__pin_sc_in_0_(grid_io_bottom_8__1__undriven_top_width_0_height_0_subtile_15__pin_sc_in_0_),
		.top_width_0_height_0_subtile_15__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_15__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_15__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_15__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_15__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_15__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_16__pin_f2a_i_0_(cbx_2__1__4_bottom_grid_top_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_16__pin_sc_in_0_(grid_io_bottom_8__1__undriven_top_width_0_height_0_subtile_16__pin_sc_in_0_),
		.top_width_0_height_0_subtile_16__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_16__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_16__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_16__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_16__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_16__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_17__pin_f2a_i_0_(cbx_2__1__4_bottom_grid_top_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_17__pin_sc_in_0_(grid_io_bottom_8__1__undriven_top_width_0_height_0_subtile_17__pin_sc_in_0_),
		.top_width_0_height_0_subtile_17__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_17__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_17__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_17__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_17__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_17__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_18__pin_f2a_i_0_(cbx_2__1__4_bottom_grid_top_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_18__pin_sc_in_0_(grid_io_bottom_8__1__undriven_top_width_0_height_0_subtile_18__pin_sc_in_0_),
		.top_width_0_height_0_subtile_18__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_18__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_18__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_18__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_18__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_18__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_19__pin_f2a_i_0_(cbx_2__1__4_bottom_grid_top_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_19__pin_sc_in_0_(grid_io_bottom_8__1__undriven_top_width_0_height_0_subtile_19__pin_sc_in_0_),
		.top_width_0_height_0_subtile_19__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_19__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_19__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_19__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_19__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_19__pin_clk_3_(clk[3]),
		.ccff_head(sb_2__0__6_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_0__pin_sc_out_0_(grid_io_bottom_8__1__undriven_top_width_0_height_0_subtile_0__pin_sc_out_0_),
		.top_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_1__pin_sc_out_0_(grid_io_bottom_8__1__undriven_top_width_0_height_0_subtile_1__pin_sc_out_0_),
		.top_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_2__pin_sc_out_0_(grid_io_bottom_8__1__undriven_top_width_0_height_0_subtile_2__pin_sc_out_0_),
		.top_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_3__pin_sc_out_0_(grid_io_bottom_8__1__undriven_top_width_0_height_0_subtile_3__pin_sc_out_0_),
		.top_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_4__pin_sc_out_0_(grid_io_bottom_8__1__undriven_top_width_0_height_0_subtile_4__pin_sc_out_0_),
		.top_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_5__pin_sc_out_0_(grid_io_bottom_8__1__undriven_top_width_0_height_0_subtile_5__pin_sc_out_0_),
		.top_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_6__pin_sc_out_0_(grid_io_bottom_8__1__undriven_top_width_0_height_0_subtile_6__pin_sc_out_0_),
		.top_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_7__pin_sc_out_0_(grid_io_bottom_8__1__undriven_top_width_0_height_0_subtile_7__pin_sc_out_0_),
		.top_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_8__pin_sc_out_0_(grid_io_bottom_8__1__undriven_top_width_0_height_0_subtile_8__pin_sc_out_0_),
		.top_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_9__pin_sc_out_0_(grid_io_bottom_8__1__undriven_top_width_0_height_0_subtile_9__pin_sc_out_0_),
		.top_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_10__pin_sc_out_0_(grid_io_bottom_8__1__undriven_top_width_0_height_0_subtile_10__pin_sc_out_0_),
		.top_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_11__pin_sc_out_0_(grid_io_bottom_8__1__undriven_top_width_0_height_0_subtile_11__pin_sc_out_0_),
		.top_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_12__pin_sc_out_0_(grid_io_bottom_8__1__undriven_top_width_0_height_0_subtile_12__pin_sc_out_0_),
		.top_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_13__pin_sc_out_0_(grid_io_bottom_8__1__undriven_top_width_0_height_0_subtile_13__pin_sc_out_0_),
		.top_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_14__pin_sc_out_0_(grid_io_bottom_8__1__undriven_top_width_0_height_0_subtile_14__pin_sc_out_0_),
		.top_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_15__pin_sc_out_0_(grid_io_bottom_8__1__undriven_top_width_0_height_0_subtile_15__pin_sc_out_0_),
		.top_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_16__pin_sc_out_0_(grid_io_bottom_8__1__undriven_top_width_0_height_0_subtile_16__pin_sc_out_0_),
		.top_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_17__pin_sc_out_0_(grid_io_bottom_8__1__undriven_top_width_0_height_0_subtile_17__pin_sc_out_0_),
		.top_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_18__pin_sc_out_0_(grid_io_bottom_8__1__undriven_top_width_0_height_0_subtile_18__pin_sc_out_0_),
		.top_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_19__pin_sc_out_0_(grid_io_bottom_8__1__undriven_top_width_0_height_0_subtile_19__pin_sc_out_0_),
		.ccff_tail(grid_io_bottom_6_ccff_tail));

	grid_io_bottom grid_io_bottom_9__1_ (
		.test_en(test_en),
		.scan_mode(scan_mode),
		.scan_clk(scan_clk),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.CFG_DONE(CFG_DONE),
		.gfpga_pad_QL_PREIO_A2F(gfpga_pad_QL_PREIO_A2F[480:499]),
		.gfpga_pad_QL_PREIO_F2A(gfpga_pad_QL_PREIO_F2A[480:499]),
		.gfpga_pad_QL_PREIO_F2A_DEF0(gfpga_pad_QL_PREIO_F2A_DEF0[480:499]),
		.gfpga_pad_QL_PREIO_F2A_DEF1(gfpga_pad_QL_PREIO_F2A_DEF1[480:499]),
		.gfpga_pad_QL_PREIO_F2A_CLK(gfpga_pad_QL_PREIO_F2A_CLK[480:499]),
		.top_width_0_height_0_subtile_0__pin_f2a_i_0_(cbx_2__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_io_bottom_9__1__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
		.top_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_1__pin_f2a_i_0_(cbx_2__1__5_bottom_grid_top_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_1__pin_sc_in_0_(grid_io_bottom_9__1__undriven_top_width_0_height_0_subtile_1__pin_sc_in_0_),
		.top_width_0_height_0_subtile_1__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_1__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_1__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_1__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_1__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_1__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_2__pin_f2a_i_0_(cbx_2__1__5_bottom_grid_top_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_2__pin_sc_in_0_(grid_io_bottom_9__1__undriven_top_width_0_height_0_subtile_2__pin_sc_in_0_),
		.top_width_0_height_0_subtile_2__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_2__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_2__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_2__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_2__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_2__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_3__pin_f2a_i_0_(cbx_2__1__5_bottom_grid_top_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_3__pin_sc_in_0_(grid_io_bottom_9__1__undriven_top_width_0_height_0_subtile_3__pin_sc_in_0_),
		.top_width_0_height_0_subtile_3__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_3__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_3__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_3__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_3__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_3__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_4__pin_f2a_i_0_(cbx_2__1__5_bottom_grid_top_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_4__pin_sc_in_0_(grid_io_bottom_9__1__undriven_top_width_0_height_0_subtile_4__pin_sc_in_0_),
		.top_width_0_height_0_subtile_4__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_4__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_4__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_4__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_4__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_4__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_5__pin_f2a_i_0_(cbx_2__1__5_bottom_grid_top_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_5__pin_sc_in_0_(grid_io_bottom_9__1__undriven_top_width_0_height_0_subtile_5__pin_sc_in_0_),
		.top_width_0_height_0_subtile_5__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_5__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_5__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_5__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_5__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_5__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_6__pin_f2a_i_0_(cbx_2__1__5_bottom_grid_top_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_6__pin_sc_in_0_(grid_io_bottom_9__1__undriven_top_width_0_height_0_subtile_6__pin_sc_in_0_),
		.top_width_0_height_0_subtile_6__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_6__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_6__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_6__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_6__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_6__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_7__pin_f2a_i_0_(cbx_2__1__5_bottom_grid_top_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_7__pin_sc_in_0_(grid_io_bottom_9__1__undriven_top_width_0_height_0_subtile_7__pin_sc_in_0_),
		.top_width_0_height_0_subtile_7__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_7__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_7__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_7__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_7__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_7__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_8__pin_f2a_i_0_(cbx_2__1__5_bottom_grid_top_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_8__pin_sc_in_0_(grid_io_bottom_9__1__undriven_top_width_0_height_0_subtile_8__pin_sc_in_0_),
		.top_width_0_height_0_subtile_8__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_8__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_8__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_8__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_8__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_8__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_9__pin_f2a_i_0_(cbx_2__1__5_bottom_grid_top_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_9__pin_sc_in_0_(grid_io_bottom_9__1__undriven_top_width_0_height_0_subtile_9__pin_sc_in_0_),
		.top_width_0_height_0_subtile_9__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_9__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_9__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_9__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_9__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_9__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_10__pin_f2a_i_0_(cbx_2__1__5_bottom_grid_top_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_10__pin_sc_in_0_(grid_io_bottom_9__1__undriven_top_width_0_height_0_subtile_10__pin_sc_in_0_),
		.top_width_0_height_0_subtile_10__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_10__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_10__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_10__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_10__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_10__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_11__pin_f2a_i_0_(cbx_2__1__5_bottom_grid_top_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_11__pin_sc_in_0_(grid_io_bottom_9__1__undriven_top_width_0_height_0_subtile_11__pin_sc_in_0_),
		.top_width_0_height_0_subtile_11__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_11__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_11__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_11__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_11__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_11__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_12__pin_f2a_i_0_(cbx_2__1__5_bottom_grid_top_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_12__pin_sc_in_0_(grid_io_bottom_9__1__undriven_top_width_0_height_0_subtile_12__pin_sc_in_0_),
		.top_width_0_height_0_subtile_12__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_12__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_12__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_12__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_12__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_12__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_13__pin_f2a_i_0_(cbx_2__1__5_bottom_grid_top_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_13__pin_sc_in_0_(grid_io_bottom_9__1__undriven_top_width_0_height_0_subtile_13__pin_sc_in_0_),
		.top_width_0_height_0_subtile_13__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_13__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_13__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_13__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_13__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_13__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_14__pin_f2a_i_0_(cbx_2__1__5_bottom_grid_top_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_14__pin_sc_in_0_(grid_io_bottom_9__1__undriven_top_width_0_height_0_subtile_14__pin_sc_in_0_),
		.top_width_0_height_0_subtile_14__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_14__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_14__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_14__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_14__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_14__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_15__pin_f2a_i_0_(cbx_2__1__5_bottom_grid_top_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_15__pin_sc_in_0_(grid_io_bottom_9__1__undriven_top_width_0_height_0_subtile_15__pin_sc_in_0_),
		.top_width_0_height_0_subtile_15__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_15__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_15__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_15__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_15__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_15__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_16__pin_f2a_i_0_(cbx_2__1__5_bottom_grid_top_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_16__pin_sc_in_0_(grid_io_bottom_9__1__undriven_top_width_0_height_0_subtile_16__pin_sc_in_0_),
		.top_width_0_height_0_subtile_16__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_16__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_16__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_16__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_16__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_16__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_17__pin_f2a_i_0_(cbx_2__1__5_bottom_grid_top_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_17__pin_sc_in_0_(grid_io_bottom_9__1__undriven_top_width_0_height_0_subtile_17__pin_sc_in_0_),
		.top_width_0_height_0_subtile_17__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_17__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_17__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_17__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_17__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_17__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_18__pin_f2a_i_0_(cbx_2__1__5_bottom_grid_top_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_18__pin_sc_in_0_(grid_io_bottom_9__1__undriven_top_width_0_height_0_subtile_18__pin_sc_in_0_),
		.top_width_0_height_0_subtile_18__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_18__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_18__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_18__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_18__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_18__pin_clk_3_(clk[3]),
		.top_width_0_height_0_subtile_19__pin_f2a_i_0_(cbx_2__1__5_bottom_grid_top_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.top_width_0_height_0_subtile_19__pin_sc_in_0_(grid_io_bottom_9__1__undriven_top_width_0_height_0_subtile_19__pin_sc_in_0_),
		.top_width_0_height_0_subtile_19__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_19__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_19__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_19__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_19__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_19__pin_clk_3_(clk[3]),
		.ccff_head(cby_9__1__0_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_0__pin_sc_out_0_(grid_io_bottom_9__1__undriven_top_width_0_height_0_subtile_0__pin_sc_out_0_),
		.top_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_1__pin_sc_out_0_(grid_io_bottom_9__1__undriven_top_width_0_height_0_subtile_1__pin_sc_out_0_),
		.top_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_2__pin_sc_out_0_(grid_io_bottom_9__1__undriven_top_width_0_height_0_subtile_2__pin_sc_out_0_),
		.top_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_3__pin_sc_out_0_(grid_io_bottom_9__1__undriven_top_width_0_height_0_subtile_3__pin_sc_out_0_),
		.top_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_4__pin_sc_out_0_(grid_io_bottom_9__1__undriven_top_width_0_height_0_subtile_4__pin_sc_out_0_),
		.top_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_5__pin_sc_out_0_(grid_io_bottom_9__1__undriven_top_width_0_height_0_subtile_5__pin_sc_out_0_),
		.top_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_6__pin_sc_out_0_(grid_io_bottom_9__1__undriven_top_width_0_height_0_subtile_6__pin_sc_out_0_),
		.top_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_7__pin_sc_out_0_(grid_io_bottom_9__1__undriven_top_width_0_height_0_subtile_7__pin_sc_out_0_),
		.top_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_8__pin_sc_out_0_(grid_io_bottom_9__1__undriven_top_width_0_height_0_subtile_8__pin_sc_out_0_),
		.top_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_9__pin_sc_out_0_(grid_io_bottom_9__1__undriven_top_width_0_height_0_subtile_9__pin_sc_out_0_),
		.top_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_10__pin_sc_out_0_(grid_io_bottom_9__1__undriven_top_width_0_height_0_subtile_10__pin_sc_out_0_),
		.top_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_11__pin_sc_out_0_(grid_io_bottom_9__1__undriven_top_width_0_height_0_subtile_11__pin_sc_out_0_),
		.top_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_12__pin_sc_out_0_(grid_io_bottom_9__1__undriven_top_width_0_height_0_subtile_12__pin_sc_out_0_),
		.top_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_13__pin_sc_out_0_(grid_io_bottom_9__1__undriven_top_width_0_height_0_subtile_13__pin_sc_out_0_),
		.top_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_14__pin_sc_out_0_(grid_io_bottom_9__1__undriven_top_width_0_height_0_subtile_14__pin_sc_out_0_),
		.top_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_15__pin_sc_out_0_(grid_io_bottom_9__1__undriven_top_width_0_height_0_subtile_15__pin_sc_out_0_),
		.top_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_16__pin_sc_out_0_(grid_io_bottom_9__1__undriven_top_width_0_height_0_subtile_16__pin_sc_out_0_),
		.top_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_17__pin_sc_out_0_(grid_io_bottom_9__1__undriven_top_width_0_height_0_subtile_17__pin_sc_out_0_),
		.top_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_18__pin_sc_out_0_(grid_io_bottom_9__1__undriven_top_width_0_height_0_subtile_18__pin_sc_out_0_),
		.top_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.top_width_0_height_0_subtile_19__pin_sc_out_0_(grid_io_bottom_9__1__undriven_top_width_0_height_0_subtile_19__pin_sc_out_0_),
		.ccff_tail(grid_io_bottom_7_ccff_tail));

	grid_clb grid_clb_2__2_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_2__2__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_0_out),
		.top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__0_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__0_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__0_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__0_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__0_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__0_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.left_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.ccff_head(cby_2__2__0_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_7_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_15_),
		.right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_17_),
		.right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_18_),
		.right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_2__2__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_2__2__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_0_ccff_tail));

	grid_clb grid_clb_2__3_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_2__3__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_1_out),
		.top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__1_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__1_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__1_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__1_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__1_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__1_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.left_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.ccff_head(cby_2__2__1_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_7_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_15_),
		.right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_17_),
		.right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_18_),
		.right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_2__3__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(ccff_tail[2]));

	grid_clb grid_clb_2__4_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_2__4__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_2_out),
		.top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__2_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__2_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__2_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__2_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__2_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__2_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.left_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.ccff_head(cby_2__2__2_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_7_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_15_),
		.right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_17_),
		.right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_18_),
		.right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_2__4__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_2_ccff_tail));

	grid_clb grid_clb_2__5_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_2__5__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_3_out),
		.top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__3_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__3_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__3_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__3_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__3_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__3_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.left_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.ccff_head(cby_2__2__3_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_7_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_15_),
		.right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_17_),
		.right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_18_),
		.right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_2__5__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_3_ccff_tail));

	grid_clb grid_clb_2__6_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_2__6__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_4_out),
		.top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__4_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__4_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__4_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__4_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__4_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__4_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.left_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.ccff_head(cby_2__2__4_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_7_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_15_),
		.right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_17_),
		.right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_18_),
		.right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_2__6__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_4_ccff_tail));

	grid_clb grid_clb_2__7_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__7__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__7__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__7__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__7__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__7__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__7__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__7__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__7__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__7__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__7__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__7__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__7__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__7__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__7__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__7__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__7__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__7__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__7__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__7__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__7__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_2__7__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_2__7__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__7__0_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__5_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__5_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__5_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__5_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__5_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__5_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.left_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.ccff_head(cby_2__2__5_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_7_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_15_),
		.right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_17_),
		.right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_18_),
		.right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_2__7__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_5_ccff_tail));

	grid_clb grid_clb_3__2_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_3__2__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_5_out),
		.top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__6_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__6_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__6_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__6_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__6_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__6_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.left_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.ccff_head(cby_2__2__6_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_7_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_15_),
		.right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_17_),
		.right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_18_),
		.right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_6_ccff_tail));

	grid_clb grid_clb_3__3_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_3__3__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_6_out),
		.top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__6_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__7_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__7_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__7_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__7_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__7_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__7_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.left_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.ccff_head(cby_2__2__7_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_7_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_15_),
		.right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_17_),
		.right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_18_),
		.right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_7_ccff_tail));

	grid_clb grid_clb_3__4_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_3__4__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_7_out),
		.top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__7_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__8_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__8_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__8_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__8_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__8_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__8_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.left_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.ccff_head(cby_2__2__8_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_7_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_15_),
		.right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_17_),
		.right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_18_),
		.right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_8_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_8_ccff_tail));

	grid_clb grid_clb_3__5_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_3__5__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_8_out),
		.top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__8_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__9_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__9_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__9_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__9_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__9_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__9_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.left_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.ccff_head(cby_2__2__9_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_7_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_15_),
		.right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_17_),
		.right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_18_),
		.right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_9_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_9_ccff_tail));

	grid_clb grid_clb_3__6_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_3__6__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_9_out),
		.top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__9_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__10_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__10_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__10_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__10_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__10_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__10_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.left_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.ccff_head(cby_2__2__10_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_7_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_15_),
		.right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_17_),
		.right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_18_),
		.right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_10_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_10_ccff_tail));

	grid_clb grid_clb_3__7_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__7__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__7__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__7__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__7__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__7__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__7__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__7__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__7__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__7__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__7__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__7__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__7__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__7__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__7__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__7__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__7__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__7__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__7__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__7__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__7__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_3__7__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_3__7__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__7__1_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__11_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__11_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__11_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__11_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__11_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__11_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.left_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.ccff_head(cby_2__2__11_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_7_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_15_),
		.right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_17_),
		.right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_18_),
		.right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_11_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_11_ccff_tail));

	grid_clb grid_clb_5__2_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_5__2__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_10_out),
		.top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__10_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__12_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__12_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__12_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__12_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__12_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__12_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.left_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.ccff_head(cby_2__2__12_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_7_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_15_),
		.right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_17_),
		.right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_18_),
		.right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_12_ccff_tail));

	grid_clb grid_clb_5__3_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_5__3__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_11_out),
		.top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__11_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__13_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__13_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__13_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__13_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__13_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__13_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.left_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.ccff_head(cby_2__2__13_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_7_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_15_),
		.right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_17_),
		.right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_18_),
		.right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_13_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_13_ccff_tail));

	grid_clb grid_clb_5__4_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_5__4__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_12_out),
		.top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__12_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__14_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__14_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__14_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__14_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__14_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__14_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.left_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.ccff_head(cby_2__2__14_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_7_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_15_),
		.right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_17_),
		.right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_18_),
		.right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_14_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_14_ccff_tail));

	grid_clb grid_clb_5__5_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_5__5__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_13_out),
		.top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__13_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__15_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__15_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__15_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__15_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__15_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__15_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.left_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.ccff_head(cby_2__2__15_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_7_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_15_),
		.right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_17_),
		.right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_18_),
		.right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_15_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_15_ccff_tail));

	grid_clb grid_clb_5__6_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_5__6__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_14_out),
		.top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__14_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__16_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__16_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__16_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__16_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__16_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__16_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.left_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.ccff_head(cby_2__2__16_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_7_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_15_),
		.right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_17_),
		.right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_18_),
		.right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_16_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_16_ccff_tail));

	grid_clb grid_clb_5__7_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__7__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__7__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__7__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__7__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__7__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__7__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__7__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__7__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__7__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__7__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__7__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__7__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__7__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__7__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__7__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__7__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__7__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__7__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__7__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__7__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_5__7__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_5__7__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__7__2_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__17_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__17_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__17_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__17_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__17_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__17_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.left_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.ccff_head(cby_2__2__17_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_7_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_15_),
		.right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_17_),
		.right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_18_),
		.right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_17_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_17_ccff_tail));

	grid_clb grid_clb_6__2_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_6__2__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_15_out),
		.top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__15_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__18_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__18_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__18_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__18_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__18_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__18_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__18_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__18_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__18_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__18_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__18_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__18_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__18_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__18_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__18_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__18_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__18_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__18_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__18_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__18_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__18_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__18_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__18_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__18_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__18_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__18_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.left_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.ccff_head(ccff_head[2]),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_7_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_15_),
		.right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_17_),
		.right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_18_),
		.right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_6__2__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_6__2__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_18_ccff_tail));

	grid_clb grid_clb_6__3_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_6__3__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_16_out),
		.top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__16_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__19_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__19_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__19_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__19_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__19_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__19_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__19_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__19_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__19_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__19_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__19_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__19_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__19_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__19_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__19_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__19_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__19_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__19_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__19_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__19_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__19_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__19_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__19_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__19_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__19_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__19_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.left_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.ccff_head(cby_2__2__19_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_7_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_15_),
		.right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_17_),
		.right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_18_),
		.right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_6__3__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_19_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_19_ccff_tail));

	grid_clb grid_clb_6__4_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_6__4__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_17_out),
		.top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__17_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__20_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__20_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__20_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__20_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__20_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__20_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__20_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__20_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__20_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__20_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__20_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__20_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__20_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__20_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__20_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__20_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__20_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__20_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__20_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__20_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__20_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__20_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__20_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__20_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__20_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__20_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.left_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.ccff_head(cby_2__2__20_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_7_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_15_),
		.right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_17_),
		.right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_18_),
		.right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_6__4__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_20_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_20_ccff_tail));

	grid_clb grid_clb_6__5_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_6__5__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_18_out),
		.top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__18_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__21_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__21_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__21_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__21_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__21_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__21_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__21_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__21_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__21_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__21_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__21_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__21_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__21_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__21_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__21_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__21_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__21_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__21_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__21_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__21_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__21_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__21_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__21_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__21_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__21_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__21_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.left_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.ccff_head(ccff_head[6]),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_7_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_15_),
		.right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_17_),
		.right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_18_),
		.right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_6__5__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_21_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_21_ccff_tail));

	grid_clb grid_clb_6__6_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_6__6__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_19_out),
		.top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__19_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__22_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__22_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__22_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__22_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__22_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__22_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__22_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__22_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__22_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__22_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__22_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__22_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__22_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__22_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__22_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__22_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__22_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__22_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__22_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__22_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__22_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__22_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__22_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__22_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__22_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__22_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.left_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.ccff_head(cby_2__2__22_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_7_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_15_),
		.right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_17_),
		.right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_18_),
		.right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_6__6__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_22_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_22_ccff_tail));

	grid_clb grid_clb_6__7_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__7__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__7__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__7__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__7__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__7__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__7__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__7__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__7__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__7__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__7__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__7__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__7__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__7__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__7__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__7__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__7__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__7__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__7__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__7__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__7__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_6__7__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_6__7__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__7__3_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__23_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__23_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__23_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__23_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__23_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__23_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__23_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__23_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__23_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__23_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__23_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__23_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__23_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__23_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__23_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__23_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__23_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__23_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__23_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__23_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__23_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__23_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__23_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__23_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__23_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__23_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.left_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.ccff_head(cby_2__2__23_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_7_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_15_),
		.right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_17_),
		.right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_18_),
		.right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_23_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_23_ccff_tail));

	grid_clb grid_clb_8__2_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_8__2__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_20_out),
		.top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__20_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__24_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__24_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__24_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__24_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__24_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__24_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__24_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__24_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__24_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__24_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__24_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__24_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__24_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__24_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__24_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__24_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__24_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__24_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__24_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__24_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__24_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__24_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__24_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__24_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__24_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__24_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.left_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.ccff_head(cby_2__2__24_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_7_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_15_),
		.right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_17_),
		.right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_18_),
		.right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_8__2__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_8__2__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_24_ccff_tail));

	grid_clb grid_clb_8__3_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_8__3__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_21_out),
		.top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__21_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__25_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__25_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__25_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__25_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__25_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__25_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__25_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__25_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__25_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__25_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__25_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__25_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__25_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__25_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__25_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__25_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__25_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__25_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__25_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__25_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__25_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__25_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__25_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__25_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__25_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__25_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.left_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.ccff_head(cby_2__2__25_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_7_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_15_),
		.right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_17_),
		.right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_18_),
		.right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_8__3__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_25_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_25_ccff_tail));

	grid_clb grid_clb_8__4_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_8__4__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_22_out),
		.top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__22_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__26_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__26_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__26_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__26_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__26_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__26_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__26_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__26_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__26_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__26_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__26_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__26_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__26_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__26_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__26_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__26_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__26_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__26_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__26_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__26_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__26_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__26_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__26_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__26_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__26_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__26_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.left_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.ccff_head(cby_2__2__26_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_7_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_15_),
		.right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_17_),
		.right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_18_),
		.right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_8__4__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_26_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_26_ccff_tail));

	grid_clb grid_clb_8__5_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_8__5__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_23_out),
		.top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__23_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__27_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__27_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__27_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__27_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__27_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__27_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__27_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__27_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__27_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__27_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__27_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__27_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__27_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__27_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__27_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__27_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__27_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__27_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__27_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__27_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__27_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__27_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__27_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__27_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__27_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__27_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.left_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.ccff_head(cby_2__2__27_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_7_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_15_),
		.right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_17_),
		.right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_18_),
		.right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_8__5__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_27_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_27_ccff_tail));

	grid_clb grid_clb_8__6_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_8__6__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_24_out),
		.top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__24_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__28_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__28_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__28_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__28_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__28_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__28_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__28_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__28_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__28_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__28_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__28_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__28_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__28_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__28_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__28_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__28_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__28_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__28_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__28_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__28_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__28_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__28_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__28_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__28_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__28_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__28_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.left_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.ccff_head(cby_2__2__28_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_7_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_15_),
		.right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_17_),
		.right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_18_),
		.right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_8__6__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_28_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_28_ccff_tail));

	grid_clb grid_clb_8__7_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__7__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__7__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__7__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__7__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__7__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__7__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__7__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__7__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__7__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__7__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__7__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__7__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__7__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__7__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__7__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__7__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__7__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__7__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__7__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__7__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_8__7__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_8__7__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__7__4_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__29_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__29_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__29_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__29_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__29_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__29_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__29_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__29_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__29_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__29_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__29_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__29_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__29_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__29_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__29_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__29_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__29_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__29_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__29_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__29_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__29_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__29_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__29_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__29_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__29_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__29_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.left_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.ccff_head(cby_2__2__29_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_7_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_15_),
		.right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_17_),
		.right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_18_),
		.right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_8__7__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_29_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_29_ccff_tail));

	grid_clb grid_clb_9__2_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_9__2__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_25_out),
		.top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__25_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.right_width_0_height_0_subtile_0__pin_I2_0_(cby_9__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.right_width_0_height_0_subtile_0__pin_I2_1_(cby_9__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.right_width_0_height_0_subtile_0__pin_I2_2_(cby_9__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.right_width_0_height_0_subtile_0__pin_I2_3_(cby_9__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.right_width_0_height_0_subtile_0__pin_I2_4_(cby_9__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.right_width_0_height_0_subtile_0__pin_I2_5_(cby_9__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.right_width_0_height_0_subtile_0__pin_I2_6_(cby_9__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.right_width_0_height_0_subtile_0__pin_I2_7_(cby_9__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.right_width_0_height_0_subtile_0__pin_I2_8_(cby_9__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.right_width_0_height_0_subtile_0__pin_I2_9_(cby_9__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.right_width_0_height_0_subtile_0__pin_I3_0_(cby_9__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.right_width_0_height_0_subtile_0__pin_I3_1_(cby_9__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.right_width_0_height_0_subtile_0__pin_I3_2_(cby_9__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.right_width_0_height_0_subtile_0__pin_I3_3_(cby_9__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.right_width_0_height_0_subtile_0__pin_I3_4_(cby_9__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.right_width_0_height_0_subtile_0__pin_I3_5_(cby_9__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.right_width_0_height_0_subtile_0__pin_I3_6_(cby_9__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.right_width_0_height_0_subtile_0__pin_I3_7_(cby_9__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.right_width_0_height_0_subtile_0__pin_I3_8_(cby_9__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.right_width_0_height_0_subtile_0__pin_I3_9_(cby_9__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.right_width_0_height_0_subtile_0__pin_IS_0_(cby_9__2__0_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.right_width_0_height_0_subtile_0__pin_IS_1_(cby_9__2__0_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.right_width_0_height_0_subtile_0__pin_IS_2_(cby_9__2__0_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.right_width_0_height_0_subtile_0__pin_IS_3_(cby_9__2__0_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.right_width_0_height_0_subtile_0__pin_IS_4_(cby_9__2__0_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.right_width_0_height_0_subtile_0__pin_IS_5_(cby_9__2__0_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.left_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.ccff_head(cby_9__2__0_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_7_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_15_),
		.right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_17_),
		.right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_18_),
		.right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_9__2__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_9__2__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_30_ccff_tail));

	grid_clb grid_clb_9__3_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_9__3__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_26_out),
		.top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__26_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.right_width_0_height_0_subtile_0__pin_I2_0_(cby_9__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.right_width_0_height_0_subtile_0__pin_I2_1_(cby_9__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.right_width_0_height_0_subtile_0__pin_I2_2_(cby_9__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.right_width_0_height_0_subtile_0__pin_I2_3_(cby_9__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.right_width_0_height_0_subtile_0__pin_I2_4_(cby_9__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.right_width_0_height_0_subtile_0__pin_I2_5_(cby_9__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.right_width_0_height_0_subtile_0__pin_I2_6_(cby_9__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.right_width_0_height_0_subtile_0__pin_I2_7_(cby_9__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.right_width_0_height_0_subtile_0__pin_I2_8_(cby_9__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.right_width_0_height_0_subtile_0__pin_I2_9_(cby_9__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.right_width_0_height_0_subtile_0__pin_I3_0_(cby_9__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.right_width_0_height_0_subtile_0__pin_I3_1_(cby_9__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.right_width_0_height_0_subtile_0__pin_I3_2_(cby_9__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.right_width_0_height_0_subtile_0__pin_I3_3_(cby_9__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.right_width_0_height_0_subtile_0__pin_I3_4_(cby_9__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.right_width_0_height_0_subtile_0__pin_I3_5_(cby_9__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.right_width_0_height_0_subtile_0__pin_I3_6_(cby_9__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.right_width_0_height_0_subtile_0__pin_I3_7_(cby_9__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.right_width_0_height_0_subtile_0__pin_I3_8_(cby_9__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.right_width_0_height_0_subtile_0__pin_I3_9_(cby_9__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.right_width_0_height_0_subtile_0__pin_IS_0_(cby_9__2__1_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.right_width_0_height_0_subtile_0__pin_IS_1_(cby_9__2__1_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.right_width_0_height_0_subtile_0__pin_IS_2_(cby_9__2__1_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.right_width_0_height_0_subtile_0__pin_IS_3_(cby_9__2__1_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.right_width_0_height_0_subtile_0__pin_IS_4_(cby_9__2__1_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.right_width_0_height_0_subtile_0__pin_IS_5_(cby_9__2__1_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.left_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.ccff_head(cby_9__2__1_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_7_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_15_),
		.right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_17_),
		.right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_18_),
		.right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_9__3__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_31_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_31_ccff_tail));

	grid_clb grid_clb_9__4_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_9__4__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_27_out),
		.top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__27_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.right_width_0_height_0_subtile_0__pin_I2_0_(cby_9__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.right_width_0_height_0_subtile_0__pin_I2_1_(cby_9__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.right_width_0_height_0_subtile_0__pin_I2_2_(cby_9__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.right_width_0_height_0_subtile_0__pin_I2_3_(cby_9__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.right_width_0_height_0_subtile_0__pin_I2_4_(cby_9__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.right_width_0_height_0_subtile_0__pin_I2_5_(cby_9__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.right_width_0_height_0_subtile_0__pin_I2_6_(cby_9__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.right_width_0_height_0_subtile_0__pin_I2_7_(cby_9__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.right_width_0_height_0_subtile_0__pin_I2_8_(cby_9__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.right_width_0_height_0_subtile_0__pin_I2_9_(cby_9__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.right_width_0_height_0_subtile_0__pin_I3_0_(cby_9__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.right_width_0_height_0_subtile_0__pin_I3_1_(cby_9__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.right_width_0_height_0_subtile_0__pin_I3_2_(cby_9__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.right_width_0_height_0_subtile_0__pin_I3_3_(cby_9__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.right_width_0_height_0_subtile_0__pin_I3_4_(cby_9__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.right_width_0_height_0_subtile_0__pin_I3_5_(cby_9__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.right_width_0_height_0_subtile_0__pin_I3_6_(cby_9__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.right_width_0_height_0_subtile_0__pin_I3_7_(cby_9__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.right_width_0_height_0_subtile_0__pin_I3_8_(cby_9__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.right_width_0_height_0_subtile_0__pin_I3_9_(cby_9__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.right_width_0_height_0_subtile_0__pin_IS_0_(cby_9__2__2_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.right_width_0_height_0_subtile_0__pin_IS_1_(cby_9__2__2_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.right_width_0_height_0_subtile_0__pin_IS_2_(cby_9__2__2_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.right_width_0_height_0_subtile_0__pin_IS_3_(cby_9__2__2_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.right_width_0_height_0_subtile_0__pin_IS_4_(cby_9__2__2_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.right_width_0_height_0_subtile_0__pin_IS_5_(cby_9__2__2_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.left_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.ccff_head(cby_9__2__2_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_7_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_15_),
		.right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_17_),
		.right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_18_),
		.right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_9__4__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_32_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_32_ccff_tail));

	grid_clb grid_clb_9__5_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_9__5__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_28_out),
		.top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__28_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.right_width_0_height_0_subtile_0__pin_I2_0_(cby_9__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.right_width_0_height_0_subtile_0__pin_I2_1_(cby_9__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.right_width_0_height_0_subtile_0__pin_I2_2_(cby_9__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.right_width_0_height_0_subtile_0__pin_I2_3_(cby_9__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.right_width_0_height_0_subtile_0__pin_I2_4_(cby_9__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.right_width_0_height_0_subtile_0__pin_I2_5_(cby_9__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.right_width_0_height_0_subtile_0__pin_I2_6_(cby_9__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.right_width_0_height_0_subtile_0__pin_I2_7_(cby_9__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.right_width_0_height_0_subtile_0__pin_I2_8_(cby_9__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.right_width_0_height_0_subtile_0__pin_I2_9_(cby_9__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.right_width_0_height_0_subtile_0__pin_I3_0_(cby_9__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.right_width_0_height_0_subtile_0__pin_I3_1_(cby_9__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.right_width_0_height_0_subtile_0__pin_I3_2_(cby_9__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.right_width_0_height_0_subtile_0__pin_I3_3_(cby_9__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.right_width_0_height_0_subtile_0__pin_I3_4_(cby_9__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.right_width_0_height_0_subtile_0__pin_I3_5_(cby_9__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.right_width_0_height_0_subtile_0__pin_I3_6_(cby_9__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.right_width_0_height_0_subtile_0__pin_I3_7_(cby_9__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.right_width_0_height_0_subtile_0__pin_I3_8_(cby_9__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.right_width_0_height_0_subtile_0__pin_I3_9_(cby_9__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.right_width_0_height_0_subtile_0__pin_IS_0_(cby_9__2__3_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.right_width_0_height_0_subtile_0__pin_IS_1_(cby_9__2__3_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.right_width_0_height_0_subtile_0__pin_IS_2_(cby_9__2__3_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.right_width_0_height_0_subtile_0__pin_IS_3_(cby_9__2__3_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.right_width_0_height_0_subtile_0__pin_IS_4_(cby_9__2__3_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.right_width_0_height_0_subtile_0__pin_IS_5_(cby_9__2__3_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.left_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.ccff_head(cby_9__2__3_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_7_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_15_),
		.right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_17_),
		.right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_18_),
		.right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_9__5__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_33_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_33_ccff_tail));

	grid_clb grid_clb_9__6_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_9__6__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_29_out),
		.top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__29_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.right_width_0_height_0_subtile_0__pin_I2_0_(cby_9__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.right_width_0_height_0_subtile_0__pin_I2_1_(cby_9__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.right_width_0_height_0_subtile_0__pin_I2_2_(cby_9__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.right_width_0_height_0_subtile_0__pin_I2_3_(cby_9__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.right_width_0_height_0_subtile_0__pin_I2_4_(cby_9__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.right_width_0_height_0_subtile_0__pin_I2_5_(cby_9__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.right_width_0_height_0_subtile_0__pin_I2_6_(cby_9__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.right_width_0_height_0_subtile_0__pin_I2_7_(cby_9__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.right_width_0_height_0_subtile_0__pin_I2_8_(cby_9__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.right_width_0_height_0_subtile_0__pin_I2_9_(cby_9__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.right_width_0_height_0_subtile_0__pin_I3_0_(cby_9__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.right_width_0_height_0_subtile_0__pin_I3_1_(cby_9__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.right_width_0_height_0_subtile_0__pin_I3_2_(cby_9__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.right_width_0_height_0_subtile_0__pin_I3_3_(cby_9__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.right_width_0_height_0_subtile_0__pin_I3_4_(cby_9__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.right_width_0_height_0_subtile_0__pin_I3_5_(cby_9__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.right_width_0_height_0_subtile_0__pin_I3_6_(cby_9__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.right_width_0_height_0_subtile_0__pin_I3_7_(cby_9__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.right_width_0_height_0_subtile_0__pin_I3_8_(cby_9__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.right_width_0_height_0_subtile_0__pin_I3_9_(cby_9__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.right_width_0_height_0_subtile_0__pin_IS_0_(cby_9__2__4_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.right_width_0_height_0_subtile_0__pin_IS_1_(cby_9__2__4_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.right_width_0_height_0_subtile_0__pin_IS_2_(cby_9__2__4_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.right_width_0_height_0_subtile_0__pin_IS_3_(cby_9__2__4_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.right_width_0_height_0_subtile_0__pin_IS_4_(cby_9__2__4_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.right_width_0_height_0_subtile_0__pin_IS_5_(cby_9__2__4_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.left_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.ccff_head(cby_9__2__4_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_7_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_15_),
		.right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_17_),
		.right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_18_),
		.right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_9__6__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_34_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_34_ccff_tail));

	grid_clb grid_clb_9__7_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__7__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__7__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__7__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__7__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__7__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__7__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__7__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__7__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__7__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__7__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__7__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__7__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__7__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__7__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__7__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__7__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__7__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__7__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__7__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__7__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_9__7__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_9__7__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__7__5_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.right_width_0_height_0_subtile_0__pin_I2_0_(cby_9__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.right_width_0_height_0_subtile_0__pin_I2_1_(cby_9__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.right_width_0_height_0_subtile_0__pin_I2_2_(cby_9__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.right_width_0_height_0_subtile_0__pin_I2_3_(cby_9__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.right_width_0_height_0_subtile_0__pin_I2_4_(cby_9__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.right_width_0_height_0_subtile_0__pin_I2_5_(cby_9__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.right_width_0_height_0_subtile_0__pin_I2_6_(cby_9__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.right_width_0_height_0_subtile_0__pin_I2_7_(cby_9__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.right_width_0_height_0_subtile_0__pin_I2_8_(cby_9__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.right_width_0_height_0_subtile_0__pin_I2_9_(cby_9__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.right_width_0_height_0_subtile_0__pin_I3_0_(cby_9__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.right_width_0_height_0_subtile_0__pin_I3_1_(cby_9__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.right_width_0_height_0_subtile_0__pin_I3_2_(cby_9__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.right_width_0_height_0_subtile_0__pin_I3_3_(cby_9__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.right_width_0_height_0_subtile_0__pin_I3_4_(cby_9__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.right_width_0_height_0_subtile_0__pin_I3_5_(cby_9__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.right_width_0_height_0_subtile_0__pin_I3_6_(cby_9__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.right_width_0_height_0_subtile_0__pin_I3_7_(cby_9__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.right_width_0_height_0_subtile_0__pin_I3_8_(cby_9__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.right_width_0_height_0_subtile_0__pin_I3_9_(cby_9__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.right_width_0_height_0_subtile_0__pin_IS_0_(cby_9__2__5_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.right_width_0_height_0_subtile_0__pin_IS_1_(cby_9__2__5_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.right_width_0_height_0_subtile_0__pin_IS_2_(cby_9__2__5_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.right_width_0_height_0_subtile_0__pin_IS_3_(cby_9__2__5_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.right_width_0_height_0_subtile_0__pin_IS_4_(cby_9__2__5_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.right_width_0_height_0_subtile_0__pin_IS_5_(cby_9__2__5_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.left_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.ccff_head(cby_9__2__5_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_7_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_8_),
		.top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_15_),
		.right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_16_),
		.right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_17_),
		.right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_18_),
		.right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_9__7__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_35_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_35_ccff_tail));

	grid_io_top grid_io_top_2__8_ (
		.test_en(test_en),
		.scan_mode(scan_mode),
		.scan_clk(scan_clk),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.CFG_DONE(CFG_DONE),
		.gfpga_pad_QL_PREIO_A2F(gfpga_pad_QL_PREIO_A2F[160:179]),
		.gfpga_pad_QL_PREIO_F2A(gfpga_pad_QL_PREIO_F2A[160:179]),
		.gfpga_pad_QL_PREIO_F2A_DEF0(gfpga_pad_QL_PREIO_F2A_DEF0[160:179]),
		.gfpga_pad_QL_PREIO_F2A_DEF1(gfpga_pad_QL_PREIO_F2A_DEF1[160:179]),
		.gfpga_pad_QL_PREIO_F2A_CLK(gfpga_pad_QL_PREIO_F2A_CLK[160:179]),
		.bottom_width_0_height_0_subtile_0__pin_f2a_i_0_(cbx_2__7__0_top_grid_bottom_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_in_0_(grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_0__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_1__pin_f2a_i_0_(cbx_2__7__0_top_grid_bottom_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_1__pin_sc_in_0_(grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_1__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_1__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_1__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_1__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_1__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_1__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_1__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_2__pin_f2a_i_0_(cbx_2__7__0_top_grid_bottom_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_2__pin_sc_in_0_(grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_2__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_2__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_2__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_2__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_2__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_2__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_2__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_3__pin_f2a_i_0_(cbx_2__7__0_top_grid_bottom_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_3__pin_sc_in_0_(grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_3__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_3__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_3__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_3__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_3__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_3__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_3__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_4__pin_f2a_i_0_(cbx_2__7__0_top_grid_bottom_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_4__pin_sc_in_0_(grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_4__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_4__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_4__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_4__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_4__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_4__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_4__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_5__pin_f2a_i_0_(cbx_2__7__0_top_grid_bottom_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_5__pin_sc_in_0_(grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_5__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_5__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_5__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_5__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_5__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_5__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_5__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_6__pin_f2a_i_0_(cbx_2__7__0_top_grid_bottom_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_6__pin_sc_in_0_(grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_6__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_6__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_6__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_6__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_6__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_6__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_6__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_7__pin_f2a_i_0_(cbx_2__7__0_top_grid_bottom_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_7__pin_sc_in_0_(grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_7__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_7__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_7__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_7__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_7__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_7__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_7__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_8__pin_f2a_i_0_(cbx_2__7__0_top_grid_bottom_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_8__pin_sc_in_0_(grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_8__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_8__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_8__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_8__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_8__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_8__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_8__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_9__pin_f2a_i_0_(cbx_2__7__0_top_grid_bottom_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_9__pin_sc_in_0_(grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_9__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_9__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_9__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_9__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_9__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_9__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_9__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_10__pin_f2a_i_0_(cbx_2__7__0_top_grid_bottom_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_10__pin_sc_in_0_(grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_10__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_10__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_10__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_10__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_10__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_10__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_10__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_11__pin_f2a_i_0_(cbx_2__7__0_top_grid_bottom_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_11__pin_sc_in_0_(grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_11__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_11__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_11__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_11__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_11__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_11__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_11__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_12__pin_f2a_i_0_(cbx_2__7__0_top_grid_bottom_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_12__pin_sc_in_0_(grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_12__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_12__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_12__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_12__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_12__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_12__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_12__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_13__pin_f2a_i_0_(cbx_2__7__0_top_grid_bottom_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_13__pin_sc_in_0_(grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_13__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_13__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_13__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_13__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_13__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_13__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_13__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_14__pin_f2a_i_0_(cbx_2__7__0_top_grid_bottom_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_14__pin_sc_in_0_(grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_14__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_14__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_14__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_14__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_14__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_14__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_14__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_15__pin_f2a_i_0_(cbx_2__7__0_top_grid_bottom_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_15__pin_sc_in_0_(grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_15__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_15__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_15__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_15__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_15__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_15__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_15__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_16__pin_f2a_i_0_(cbx_2__7__0_top_grid_bottom_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_16__pin_sc_in_0_(grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_16__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_16__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_16__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_16__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_16__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_16__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_16__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_17__pin_f2a_i_0_(cbx_2__7__0_top_grid_bottom_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_17__pin_sc_in_0_(grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_17__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_17__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_17__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_17__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_17__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_17__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_17__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_18__pin_f2a_i_0_(cbx_2__7__0_top_grid_bottom_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_18__pin_sc_in_0_(grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_18__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_18__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_18__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_18__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_18__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_18__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_18__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_19__pin_f2a_i_0_(cbx_2__7__0_top_grid_bottom_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_19__pin_sc_in_0_(grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_19__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_19__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_19__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_19__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_19__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_19__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_19__pin_clk_3_(clk[3]),
		.ccff_head(cbx_2__7__0_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_1__pin_sc_out_0_(grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_1__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_2__pin_sc_out_0_(grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_2__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_3__pin_sc_out_0_(grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_3__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_4__pin_sc_out_0_(grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_4__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_5__pin_sc_out_0_(grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_5__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_6__pin_sc_out_0_(grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_6__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_7__pin_sc_out_0_(grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_7__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_8__pin_sc_out_0_(grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_8__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_9__pin_sc_out_0_(grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_9__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_10__pin_sc_out_0_(grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_10__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_11__pin_sc_out_0_(grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_11__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_12__pin_sc_out_0_(grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_12__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_13__pin_sc_out_0_(grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_13__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_14__pin_sc_out_0_(grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_14__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_15__pin_sc_out_0_(grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_15__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_16__pin_sc_out_0_(grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_16__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_17__pin_sc_out_0_(grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_17__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_18__pin_sc_out_0_(grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_18__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_19__pin_sc_out_0_(grid_io_top_2__8__undriven_bottom_width_0_height_0_subtile_19__pin_sc_out_0_),
		.ccff_tail(grid_io_top_0_ccff_tail));

	grid_io_top grid_io_top_3__8_ (
		.test_en(test_en),
		.scan_mode(scan_mode),
		.scan_clk(scan_clk),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.CFG_DONE(CFG_DONE),
		.gfpga_pad_QL_PREIO_A2F(gfpga_pad_QL_PREIO_A2F[180:199]),
		.gfpga_pad_QL_PREIO_F2A(gfpga_pad_QL_PREIO_F2A[180:199]),
		.gfpga_pad_QL_PREIO_F2A_DEF0(gfpga_pad_QL_PREIO_F2A_DEF0[180:199]),
		.gfpga_pad_QL_PREIO_F2A_DEF1(gfpga_pad_QL_PREIO_F2A_DEF1[180:199]),
		.gfpga_pad_QL_PREIO_F2A_CLK(gfpga_pad_QL_PREIO_F2A_CLK[180:199]),
		.bottom_width_0_height_0_subtile_0__pin_f2a_i_0_(cbx_2__7__1_top_grid_bottom_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_in_0_(grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_0__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_1__pin_f2a_i_0_(cbx_2__7__1_top_grid_bottom_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_1__pin_sc_in_0_(grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_1__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_1__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_1__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_1__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_1__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_1__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_1__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_2__pin_f2a_i_0_(cbx_2__7__1_top_grid_bottom_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_2__pin_sc_in_0_(grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_2__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_2__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_2__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_2__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_2__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_2__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_2__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_3__pin_f2a_i_0_(cbx_2__7__1_top_grid_bottom_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_3__pin_sc_in_0_(grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_3__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_3__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_3__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_3__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_3__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_3__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_3__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_4__pin_f2a_i_0_(cbx_2__7__1_top_grid_bottom_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_4__pin_sc_in_0_(grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_4__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_4__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_4__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_4__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_4__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_4__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_4__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_5__pin_f2a_i_0_(cbx_2__7__1_top_grid_bottom_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_5__pin_sc_in_0_(grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_5__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_5__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_5__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_5__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_5__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_5__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_5__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_6__pin_f2a_i_0_(cbx_2__7__1_top_grid_bottom_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_6__pin_sc_in_0_(grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_6__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_6__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_6__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_6__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_6__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_6__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_6__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_7__pin_f2a_i_0_(cbx_2__7__1_top_grid_bottom_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_7__pin_sc_in_0_(grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_7__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_7__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_7__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_7__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_7__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_7__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_7__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_8__pin_f2a_i_0_(cbx_2__7__1_top_grid_bottom_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_8__pin_sc_in_0_(grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_8__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_8__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_8__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_8__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_8__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_8__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_8__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_9__pin_f2a_i_0_(cbx_2__7__1_top_grid_bottom_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_9__pin_sc_in_0_(grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_9__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_9__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_9__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_9__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_9__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_9__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_9__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_10__pin_f2a_i_0_(cbx_2__7__1_top_grid_bottom_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_10__pin_sc_in_0_(grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_10__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_10__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_10__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_10__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_10__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_10__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_10__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_11__pin_f2a_i_0_(cbx_2__7__1_top_grid_bottom_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_11__pin_sc_in_0_(grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_11__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_11__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_11__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_11__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_11__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_11__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_11__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_12__pin_f2a_i_0_(cbx_2__7__1_top_grid_bottom_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_12__pin_sc_in_0_(grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_12__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_12__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_12__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_12__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_12__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_12__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_12__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_13__pin_f2a_i_0_(cbx_2__7__1_top_grid_bottom_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_13__pin_sc_in_0_(grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_13__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_13__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_13__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_13__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_13__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_13__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_13__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_14__pin_f2a_i_0_(cbx_2__7__1_top_grid_bottom_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_14__pin_sc_in_0_(grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_14__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_14__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_14__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_14__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_14__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_14__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_14__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_15__pin_f2a_i_0_(cbx_2__7__1_top_grid_bottom_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_15__pin_sc_in_0_(grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_15__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_15__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_15__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_15__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_15__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_15__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_15__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_16__pin_f2a_i_0_(cbx_2__7__1_top_grid_bottom_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_16__pin_sc_in_0_(grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_16__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_16__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_16__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_16__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_16__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_16__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_16__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_17__pin_f2a_i_0_(cbx_2__7__1_top_grid_bottom_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_17__pin_sc_in_0_(grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_17__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_17__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_17__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_17__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_17__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_17__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_17__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_18__pin_f2a_i_0_(cbx_2__7__1_top_grid_bottom_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_18__pin_sc_in_0_(grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_18__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_18__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_18__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_18__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_18__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_18__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_18__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_19__pin_f2a_i_0_(cbx_2__7__1_top_grid_bottom_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_19__pin_sc_in_0_(grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_19__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_19__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_19__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_19__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_19__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_19__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_19__pin_clk_3_(clk[3]),
		.ccff_head(cbx_2__7__1_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_1__pin_sc_out_0_(grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_1__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_2__pin_sc_out_0_(grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_2__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_3__pin_sc_out_0_(grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_3__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_4__pin_sc_out_0_(grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_4__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_5__pin_sc_out_0_(grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_5__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_6__pin_sc_out_0_(grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_6__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_7__pin_sc_out_0_(grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_7__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_8__pin_sc_out_0_(grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_8__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_9__pin_sc_out_0_(grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_9__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_10__pin_sc_out_0_(grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_10__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_11__pin_sc_out_0_(grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_11__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_12__pin_sc_out_0_(grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_12__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_13__pin_sc_out_0_(grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_13__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_14__pin_sc_out_0_(grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_14__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_15__pin_sc_out_0_(grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_15__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_16__pin_sc_out_0_(grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_16__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_17__pin_sc_out_0_(grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_17__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_18__pin_sc_out_0_(grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_18__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_19__pin_sc_out_0_(grid_io_top_3__8__undriven_bottom_width_0_height_0_subtile_19__pin_sc_out_0_),
		.ccff_tail(grid_io_top_1_ccff_tail));

	grid_io_top grid_io_top_4__8_ (
		.test_en(test_en),
		.scan_mode(scan_mode),
		.scan_clk(scan_clk),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.CFG_DONE(CFG_DONE),
		.gfpga_pad_QL_PREIO_A2F(gfpga_pad_QL_PREIO_A2F[200:219]),
		.gfpga_pad_QL_PREIO_F2A(gfpga_pad_QL_PREIO_F2A[200:219]),
		.gfpga_pad_QL_PREIO_F2A_DEF0(gfpga_pad_QL_PREIO_F2A_DEF0[200:219]),
		.gfpga_pad_QL_PREIO_F2A_DEF1(gfpga_pad_QL_PREIO_F2A_DEF1[200:219]),
		.gfpga_pad_QL_PREIO_F2A_CLK(gfpga_pad_QL_PREIO_F2A_CLK[200:219]),
		.bottom_width_0_height_0_subtile_0__pin_f2a_i_0_(cbx_4__7__0_top_grid_bottom_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_in_0_(grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_0__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_1__pin_f2a_i_0_(cbx_4__7__0_top_grid_bottom_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_1__pin_sc_in_0_(grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_1__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_1__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_1__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_1__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_1__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_1__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_1__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_2__pin_f2a_i_0_(cbx_4__7__0_top_grid_bottom_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_2__pin_sc_in_0_(grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_2__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_2__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_2__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_2__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_2__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_2__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_2__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_3__pin_f2a_i_0_(cbx_4__7__0_top_grid_bottom_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_3__pin_sc_in_0_(grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_3__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_3__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_3__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_3__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_3__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_3__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_3__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_4__pin_f2a_i_0_(cbx_4__7__0_top_grid_bottom_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_4__pin_sc_in_0_(grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_4__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_4__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_4__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_4__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_4__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_4__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_4__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_5__pin_f2a_i_0_(cbx_4__7__0_top_grid_bottom_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_5__pin_sc_in_0_(grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_5__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_5__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_5__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_5__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_5__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_5__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_5__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_6__pin_f2a_i_0_(cbx_4__7__0_top_grid_bottom_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_6__pin_sc_in_0_(grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_6__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_6__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_6__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_6__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_6__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_6__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_6__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_7__pin_f2a_i_0_(cbx_4__7__0_top_grid_bottom_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_7__pin_sc_in_0_(grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_7__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_7__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_7__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_7__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_7__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_7__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_7__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_8__pin_f2a_i_0_(cbx_4__7__0_top_grid_bottom_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_8__pin_sc_in_0_(grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_8__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_8__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_8__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_8__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_8__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_8__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_8__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_9__pin_f2a_i_0_(cbx_4__7__0_top_grid_bottom_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_9__pin_sc_in_0_(grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_9__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_9__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_9__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_9__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_9__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_9__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_9__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_10__pin_f2a_i_0_(cbx_4__7__0_top_grid_bottom_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_10__pin_sc_in_0_(grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_10__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_10__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_10__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_10__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_10__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_10__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_10__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_11__pin_f2a_i_0_(cbx_4__7__0_top_grid_bottom_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_11__pin_sc_in_0_(grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_11__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_11__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_11__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_11__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_11__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_11__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_11__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_12__pin_f2a_i_0_(cbx_4__7__0_top_grid_bottom_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_12__pin_sc_in_0_(grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_12__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_12__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_12__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_12__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_12__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_12__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_12__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_13__pin_f2a_i_0_(cbx_4__7__0_top_grid_bottom_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_13__pin_sc_in_0_(grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_13__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_13__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_13__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_13__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_13__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_13__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_13__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_14__pin_f2a_i_0_(cbx_4__7__0_top_grid_bottom_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_14__pin_sc_in_0_(grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_14__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_14__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_14__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_14__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_14__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_14__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_14__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_15__pin_f2a_i_0_(cbx_4__7__0_top_grid_bottom_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_15__pin_sc_in_0_(grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_15__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_15__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_15__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_15__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_15__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_15__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_15__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_16__pin_f2a_i_0_(cbx_4__7__0_top_grid_bottom_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_16__pin_sc_in_0_(grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_16__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_16__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_16__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_16__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_16__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_16__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_16__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_17__pin_f2a_i_0_(cbx_4__7__0_top_grid_bottom_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_17__pin_sc_in_0_(grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_17__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_17__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_17__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_17__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_17__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_17__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_17__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_18__pin_f2a_i_0_(cbx_4__7__0_top_grid_bottom_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_18__pin_sc_in_0_(grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_18__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_18__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_18__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_18__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_18__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_18__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_18__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_19__pin_f2a_i_0_(cbx_4__7__0_top_grid_bottom_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_19__pin_sc_in_0_(grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_19__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_19__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_19__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_19__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_19__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_19__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_19__pin_clk_3_(clk[3]),
		.ccff_head(cbx_4__7__0_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_1__pin_sc_out_0_(grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_1__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_2__pin_sc_out_0_(grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_2__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_3__pin_sc_out_0_(grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_3__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_4__pin_sc_out_0_(grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_4__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_5__pin_sc_out_0_(grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_5__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_6__pin_sc_out_0_(grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_6__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_7__pin_sc_out_0_(grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_7__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_8__pin_sc_out_0_(grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_8__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_9__pin_sc_out_0_(grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_9__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_10__pin_sc_out_0_(grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_10__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_11__pin_sc_out_0_(grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_11__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_12__pin_sc_out_0_(grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_12__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_13__pin_sc_out_0_(grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_13__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_14__pin_sc_out_0_(grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_14__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_15__pin_sc_out_0_(grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_15__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_16__pin_sc_out_0_(grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_16__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_17__pin_sc_out_0_(grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_17__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_18__pin_sc_out_0_(grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_18__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_19__pin_sc_out_0_(grid_io_top_4__8__undriven_bottom_width_0_height_0_subtile_19__pin_sc_out_0_),
		.ccff_tail(grid_io_top_2_ccff_tail));

	grid_io_top grid_io_top_5__8_ (
		.test_en(test_en),
		.scan_mode(scan_mode),
		.scan_clk(scan_clk),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.CFG_DONE(CFG_DONE),
		.gfpga_pad_QL_PREIO_A2F(gfpga_pad_QL_PREIO_A2F[220:239]),
		.gfpga_pad_QL_PREIO_F2A(gfpga_pad_QL_PREIO_F2A[220:239]),
		.gfpga_pad_QL_PREIO_F2A_DEF0(gfpga_pad_QL_PREIO_F2A_DEF0[220:239]),
		.gfpga_pad_QL_PREIO_F2A_DEF1(gfpga_pad_QL_PREIO_F2A_DEF1[220:239]),
		.gfpga_pad_QL_PREIO_F2A_CLK(gfpga_pad_QL_PREIO_F2A_CLK[220:239]),
		.bottom_width_0_height_0_subtile_0__pin_f2a_i_0_(cbx_2__7__2_top_grid_bottom_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_in_0_(grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_0__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_1__pin_f2a_i_0_(cbx_2__7__2_top_grid_bottom_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_1__pin_sc_in_0_(grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_1__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_1__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_1__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_1__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_1__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_1__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_1__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_2__pin_f2a_i_0_(cbx_2__7__2_top_grid_bottom_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_2__pin_sc_in_0_(grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_2__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_2__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_2__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_2__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_2__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_2__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_2__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_3__pin_f2a_i_0_(cbx_2__7__2_top_grid_bottom_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_3__pin_sc_in_0_(grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_3__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_3__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_3__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_3__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_3__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_3__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_3__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_4__pin_f2a_i_0_(cbx_2__7__2_top_grid_bottom_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_4__pin_sc_in_0_(grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_4__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_4__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_4__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_4__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_4__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_4__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_4__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_5__pin_f2a_i_0_(cbx_2__7__2_top_grid_bottom_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_5__pin_sc_in_0_(grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_5__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_5__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_5__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_5__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_5__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_5__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_5__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_6__pin_f2a_i_0_(cbx_2__7__2_top_grid_bottom_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_6__pin_sc_in_0_(grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_6__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_6__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_6__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_6__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_6__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_6__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_6__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_7__pin_f2a_i_0_(cbx_2__7__2_top_grid_bottom_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_7__pin_sc_in_0_(grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_7__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_7__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_7__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_7__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_7__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_7__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_7__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_8__pin_f2a_i_0_(cbx_2__7__2_top_grid_bottom_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_8__pin_sc_in_0_(grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_8__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_8__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_8__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_8__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_8__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_8__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_8__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_9__pin_f2a_i_0_(cbx_2__7__2_top_grid_bottom_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_9__pin_sc_in_0_(grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_9__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_9__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_9__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_9__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_9__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_9__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_9__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_10__pin_f2a_i_0_(cbx_2__7__2_top_grid_bottom_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_10__pin_sc_in_0_(grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_10__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_10__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_10__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_10__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_10__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_10__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_10__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_11__pin_f2a_i_0_(cbx_2__7__2_top_grid_bottom_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_11__pin_sc_in_0_(grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_11__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_11__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_11__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_11__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_11__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_11__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_11__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_12__pin_f2a_i_0_(cbx_2__7__2_top_grid_bottom_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_12__pin_sc_in_0_(grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_12__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_12__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_12__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_12__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_12__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_12__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_12__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_13__pin_f2a_i_0_(cbx_2__7__2_top_grid_bottom_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_13__pin_sc_in_0_(grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_13__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_13__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_13__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_13__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_13__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_13__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_13__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_14__pin_f2a_i_0_(cbx_2__7__2_top_grid_bottom_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_14__pin_sc_in_0_(grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_14__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_14__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_14__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_14__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_14__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_14__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_14__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_15__pin_f2a_i_0_(cbx_2__7__2_top_grid_bottom_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_15__pin_sc_in_0_(grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_15__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_15__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_15__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_15__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_15__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_15__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_15__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_16__pin_f2a_i_0_(cbx_2__7__2_top_grid_bottom_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_16__pin_sc_in_0_(grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_16__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_16__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_16__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_16__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_16__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_16__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_16__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_17__pin_f2a_i_0_(cbx_2__7__2_top_grid_bottom_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_17__pin_sc_in_0_(grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_17__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_17__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_17__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_17__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_17__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_17__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_17__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_18__pin_f2a_i_0_(cbx_2__7__2_top_grid_bottom_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_18__pin_sc_in_0_(grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_18__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_18__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_18__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_18__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_18__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_18__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_18__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_19__pin_f2a_i_0_(cbx_2__7__2_top_grid_bottom_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_19__pin_sc_in_0_(grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_19__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_19__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_19__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_19__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_19__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_19__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_19__pin_clk_3_(clk[3]),
		.ccff_head(cbx_2__7__2_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_1__pin_sc_out_0_(grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_1__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_2__pin_sc_out_0_(grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_2__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_3__pin_sc_out_0_(grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_3__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_4__pin_sc_out_0_(grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_4__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_5__pin_sc_out_0_(grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_5__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_6__pin_sc_out_0_(grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_6__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_7__pin_sc_out_0_(grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_7__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_8__pin_sc_out_0_(grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_8__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_9__pin_sc_out_0_(grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_9__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_10__pin_sc_out_0_(grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_10__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_11__pin_sc_out_0_(grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_11__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_12__pin_sc_out_0_(grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_12__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_13__pin_sc_out_0_(grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_13__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_14__pin_sc_out_0_(grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_14__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_15__pin_sc_out_0_(grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_15__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_16__pin_sc_out_0_(grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_16__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_17__pin_sc_out_0_(grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_17__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_18__pin_sc_out_0_(grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_18__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_19__pin_sc_out_0_(grid_io_top_5__8__undriven_bottom_width_0_height_0_subtile_19__pin_sc_out_0_),
		.ccff_tail(grid_io_top_3_ccff_tail));

	grid_io_top grid_io_top_6__8_ (
		.test_en(test_en),
		.scan_mode(scan_mode),
		.scan_clk(scan_clk),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.CFG_DONE(CFG_DONE),
		.gfpga_pad_QL_PREIO_A2F(gfpga_pad_QL_PREIO_A2F[240:259]),
		.gfpga_pad_QL_PREIO_F2A(gfpga_pad_QL_PREIO_F2A[240:259]),
		.gfpga_pad_QL_PREIO_F2A_DEF0(gfpga_pad_QL_PREIO_F2A_DEF0[240:259]),
		.gfpga_pad_QL_PREIO_F2A_DEF1(gfpga_pad_QL_PREIO_F2A_DEF1[240:259]),
		.gfpga_pad_QL_PREIO_F2A_CLK(gfpga_pad_QL_PREIO_F2A_CLK[240:259]),
		.bottom_width_0_height_0_subtile_0__pin_f2a_i_0_(cbx_2__7__3_top_grid_bottom_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_in_0_(grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_0__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_1__pin_f2a_i_0_(cbx_2__7__3_top_grid_bottom_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_1__pin_sc_in_0_(grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_1__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_1__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_1__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_1__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_1__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_1__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_1__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_2__pin_f2a_i_0_(cbx_2__7__3_top_grid_bottom_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_2__pin_sc_in_0_(grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_2__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_2__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_2__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_2__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_2__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_2__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_2__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_3__pin_f2a_i_0_(cbx_2__7__3_top_grid_bottom_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_3__pin_sc_in_0_(grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_3__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_3__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_3__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_3__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_3__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_3__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_3__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_4__pin_f2a_i_0_(cbx_2__7__3_top_grid_bottom_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_4__pin_sc_in_0_(grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_4__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_4__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_4__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_4__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_4__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_4__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_4__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_5__pin_f2a_i_0_(cbx_2__7__3_top_grid_bottom_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_5__pin_sc_in_0_(grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_5__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_5__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_5__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_5__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_5__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_5__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_5__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_6__pin_f2a_i_0_(cbx_2__7__3_top_grid_bottom_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_6__pin_sc_in_0_(grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_6__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_6__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_6__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_6__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_6__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_6__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_6__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_7__pin_f2a_i_0_(cbx_2__7__3_top_grid_bottom_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_7__pin_sc_in_0_(grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_7__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_7__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_7__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_7__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_7__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_7__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_7__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_8__pin_f2a_i_0_(cbx_2__7__3_top_grid_bottom_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_8__pin_sc_in_0_(grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_8__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_8__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_8__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_8__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_8__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_8__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_8__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_9__pin_f2a_i_0_(cbx_2__7__3_top_grid_bottom_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_9__pin_sc_in_0_(grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_9__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_9__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_9__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_9__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_9__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_9__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_9__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_10__pin_f2a_i_0_(cbx_2__7__3_top_grid_bottom_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_10__pin_sc_in_0_(grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_10__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_10__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_10__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_10__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_10__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_10__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_10__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_11__pin_f2a_i_0_(cbx_2__7__3_top_grid_bottom_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_11__pin_sc_in_0_(grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_11__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_11__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_11__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_11__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_11__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_11__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_11__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_12__pin_f2a_i_0_(cbx_2__7__3_top_grid_bottom_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_12__pin_sc_in_0_(grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_12__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_12__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_12__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_12__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_12__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_12__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_12__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_13__pin_f2a_i_0_(cbx_2__7__3_top_grid_bottom_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_13__pin_sc_in_0_(grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_13__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_13__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_13__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_13__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_13__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_13__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_13__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_14__pin_f2a_i_0_(cbx_2__7__3_top_grid_bottom_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_14__pin_sc_in_0_(grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_14__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_14__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_14__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_14__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_14__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_14__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_14__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_15__pin_f2a_i_0_(cbx_2__7__3_top_grid_bottom_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_15__pin_sc_in_0_(grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_15__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_15__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_15__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_15__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_15__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_15__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_15__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_16__pin_f2a_i_0_(cbx_2__7__3_top_grid_bottom_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_16__pin_sc_in_0_(grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_16__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_16__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_16__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_16__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_16__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_16__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_16__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_17__pin_f2a_i_0_(cbx_2__7__3_top_grid_bottom_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_17__pin_sc_in_0_(grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_17__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_17__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_17__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_17__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_17__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_17__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_17__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_18__pin_f2a_i_0_(cbx_2__7__3_top_grid_bottom_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_18__pin_sc_in_0_(grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_18__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_18__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_18__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_18__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_18__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_18__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_18__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_19__pin_f2a_i_0_(cbx_2__7__3_top_grid_bottom_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_19__pin_sc_in_0_(grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_19__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_19__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_19__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_19__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_19__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_19__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_19__pin_clk_3_(clk[3]),
		.ccff_head(cbx_2__7__3_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_1__pin_sc_out_0_(grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_1__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_2__pin_sc_out_0_(grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_2__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_3__pin_sc_out_0_(grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_3__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_4__pin_sc_out_0_(grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_4__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_5__pin_sc_out_0_(grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_5__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_6__pin_sc_out_0_(grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_6__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_7__pin_sc_out_0_(grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_7__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_8__pin_sc_out_0_(grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_8__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_9__pin_sc_out_0_(grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_9__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_10__pin_sc_out_0_(grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_10__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_11__pin_sc_out_0_(grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_11__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_12__pin_sc_out_0_(grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_12__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_13__pin_sc_out_0_(grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_13__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_14__pin_sc_out_0_(grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_14__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_15__pin_sc_out_0_(grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_15__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_16__pin_sc_out_0_(grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_16__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_17__pin_sc_out_0_(grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_17__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_18__pin_sc_out_0_(grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_18__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_19__pin_sc_out_0_(grid_io_top_6__8__undriven_bottom_width_0_height_0_subtile_19__pin_sc_out_0_),
		.ccff_tail(grid_io_top_4_ccff_tail));

	grid_io_top grid_io_top_7__8_ (
		.test_en(test_en),
		.scan_mode(scan_mode),
		.scan_clk(scan_clk),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.CFG_DONE(CFG_DONE),
		.gfpga_pad_QL_PREIO_A2F(gfpga_pad_QL_PREIO_A2F[260:279]),
		.gfpga_pad_QL_PREIO_F2A(gfpga_pad_QL_PREIO_F2A[260:279]),
		.gfpga_pad_QL_PREIO_F2A_DEF0(gfpga_pad_QL_PREIO_F2A_DEF0[260:279]),
		.gfpga_pad_QL_PREIO_F2A_DEF1(gfpga_pad_QL_PREIO_F2A_DEF1[260:279]),
		.gfpga_pad_QL_PREIO_F2A_CLK(gfpga_pad_QL_PREIO_F2A_CLK[260:279]),
		.bottom_width_0_height_0_subtile_0__pin_f2a_i_0_(cbx_4__7__1_top_grid_bottom_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_in_0_(grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_0__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_1__pin_f2a_i_0_(cbx_4__7__1_top_grid_bottom_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_1__pin_sc_in_0_(grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_1__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_1__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_1__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_1__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_1__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_1__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_1__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_2__pin_f2a_i_0_(cbx_4__7__1_top_grid_bottom_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_2__pin_sc_in_0_(grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_2__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_2__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_2__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_2__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_2__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_2__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_2__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_3__pin_f2a_i_0_(cbx_4__7__1_top_grid_bottom_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_3__pin_sc_in_0_(grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_3__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_3__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_3__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_3__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_3__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_3__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_3__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_4__pin_f2a_i_0_(cbx_4__7__1_top_grid_bottom_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_4__pin_sc_in_0_(grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_4__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_4__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_4__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_4__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_4__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_4__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_4__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_5__pin_f2a_i_0_(cbx_4__7__1_top_grid_bottom_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_5__pin_sc_in_0_(grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_5__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_5__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_5__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_5__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_5__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_5__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_5__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_6__pin_f2a_i_0_(cbx_4__7__1_top_grid_bottom_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_6__pin_sc_in_0_(grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_6__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_6__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_6__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_6__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_6__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_6__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_6__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_7__pin_f2a_i_0_(cbx_4__7__1_top_grid_bottom_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_7__pin_sc_in_0_(grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_7__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_7__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_7__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_7__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_7__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_7__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_7__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_8__pin_f2a_i_0_(cbx_4__7__1_top_grid_bottom_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_8__pin_sc_in_0_(grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_8__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_8__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_8__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_8__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_8__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_8__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_8__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_9__pin_f2a_i_0_(cbx_4__7__1_top_grid_bottom_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_9__pin_sc_in_0_(grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_9__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_9__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_9__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_9__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_9__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_9__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_9__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_10__pin_f2a_i_0_(cbx_4__7__1_top_grid_bottom_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_10__pin_sc_in_0_(grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_10__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_10__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_10__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_10__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_10__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_10__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_10__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_11__pin_f2a_i_0_(cbx_4__7__1_top_grid_bottom_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_11__pin_sc_in_0_(grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_11__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_11__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_11__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_11__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_11__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_11__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_11__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_12__pin_f2a_i_0_(cbx_4__7__1_top_grid_bottom_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_12__pin_sc_in_0_(grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_12__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_12__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_12__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_12__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_12__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_12__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_12__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_13__pin_f2a_i_0_(cbx_4__7__1_top_grid_bottom_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_13__pin_sc_in_0_(grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_13__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_13__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_13__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_13__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_13__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_13__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_13__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_14__pin_f2a_i_0_(cbx_4__7__1_top_grid_bottom_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_14__pin_sc_in_0_(grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_14__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_14__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_14__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_14__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_14__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_14__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_14__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_15__pin_f2a_i_0_(cbx_4__7__1_top_grid_bottom_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_15__pin_sc_in_0_(grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_15__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_15__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_15__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_15__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_15__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_15__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_15__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_16__pin_f2a_i_0_(cbx_4__7__1_top_grid_bottom_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_16__pin_sc_in_0_(grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_16__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_16__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_16__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_16__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_16__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_16__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_16__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_17__pin_f2a_i_0_(cbx_4__7__1_top_grid_bottom_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_17__pin_sc_in_0_(grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_17__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_17__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_17__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_17__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_17__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_17__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_17__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_18__pin_f2a_i_0_(cbx_4__7__1_top_grid_bottom_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_18__pin_sc_in_0_(grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_18__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_18__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_18__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_18__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_18__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_18__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_18__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_19__pin_f2a_i_0_(cbx_4__7__1_top_grid_bottom_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_19__pin_sc_in_0_(grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_19__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_19__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_19__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_19__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_19__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_19__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_19__pin_clk_3_(clk[3]),
		.ccff_head(cbx_4__7__1_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_1__pin_sc_out_0_(grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_1__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_2__pin_sc_out_0_(grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_2__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_3__pin_sc_out_0_(grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_3__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_4__pin_sc_out_0_(grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_4__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_5__pin_sc_out_0_(grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_5__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_6__pin_sc_out_0_(grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_6__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_7__pin_sc_out_0_(grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_7__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_8__pin_sc_out_0_(grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_8__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_9__pin_sc_out_0_(grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_9__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_10__pin_sc_out_0_(grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_10__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_11__pin_sc_out_0_(grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_11__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_12__pin_sc_out_0_(grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_12__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_13__pin_sc_out_0_(grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_13__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_14__pin_sc_out_0_(grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_14__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_15__pin_sc_out_0_(grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_15__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_16__pin_sc_out_0_(grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_16__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_17__pin_sc_out_0_(grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_17__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_18__pin_sc_out_0_(grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_18__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_19__pin_sc_out_0_(grid_io_top_7__8__undriven_bottom_width_0_height_0_subtile_19__pin_sc_out_0_),
		.ccff_tail(grid_io_top_5_ccff_tail));

	grid_io_top grid_io_top_8__8_ (
		.test_en(test_en),
		.scan_mode(scan_mode),
		.scan_clk(scan_clk),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.CFG_DONE(CFG_DONE),
		.gfpga_pad_QL_PREIO_A2F(gfpga_pad_QL_PREIO_A2F[280:299]),
		.gfpga_pad_QL_PREIO_F2A(gfpga_pad_QL_PREIO_F2A[280:299]),
		.gfpga_pad_QL_PREIO_F2A_DEF0(gfpga_pad_QL_PREIO_F2A_DEF0[280:299]),
		.gfpga_pad_QL_PREIO_F2A_DEF1(gfpga_pad_QL_PREIO_F2A_DEF1[280:299]),
		.gfpga_pad_QL_PREIO_F2A_CLK(gfpga_pad_QL_PREIO_F2A_CLK[280:299]),
		.bottom_width_0_height_0_subtile_0__pin_f2a_i_0_(cbx_2__7__4_top_grid_bottom_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_in_0_(grid_io_top_8__8__undriven_bottom_width_0_height_0_subtile_0__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_1__pin_f2a_i_0_(cbx_2__7__4_top_grid_bottom_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_1__pin_sc_in_0_(grid_io_top_8__8__undriven_bottom_width_0_height_0_subtile_1__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_1__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_1__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_1__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_1__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_1__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_1__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_2__pin_f2a_i_0_(cbx_2__7__4_top_grid_bottom_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_2__pin_sc_in_0_(grid_io_top_8__8__undriven_bottom_width_0_height_0_subtile_2__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_2__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_2__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_2__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_2__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_2__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_2__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_3__pin_f2a_i_0_(cbx_2__7__4_top_grid_bottom_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_3__pin_sc_in_0_(grid_io_top_8__8__undriven_bottom_width_0_height_0_subtile_3__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_3__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_3__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_3__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_3__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_3__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_3__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_4__pin_f2a_i_0_(cbx_2__7__4_top_grid_bottom_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_4__pin_sc_in_0_(grid_io_top_8__8__undriven_bottom_width_0_height_0_subtile_4__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_4__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_4__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_4__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_4__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_4__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_4__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_5__pin_f2a_i_0_(cbx_2__7__4_top_grid_bottom_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_5__pin_sc_in_0_(grid_io_top_8__8__undriven_bottom_width_0_height_0_subtile_5__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_5__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_5__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_5__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_5__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_5__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_5__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_6__pin_f2a_i_0_(cbx_2__7__4_top_grid_bottom_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_6__pin_sc_in_0_(grid_io_top_8__8__undriven_bottom_width_0_height_0_subtile_6__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_6__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_6__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_6__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_6__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_6__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_6__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_7__pin_f2a_i_0_(cbx_2__7__4_top_grid_bottom_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_7__pin_sc_in_0_(grid_io_top_8__8__undriven_bottom_width_0_height_0_subtile_7__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_7__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_7__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_7__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_7__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_7__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_7__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_8__pin_f2a_i_0_(cbx_2__7__4_top_grid_bottom_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_8__pin_sc_in_0_(grid_io_top_8__8__undriven_bottom_width_0_height_0_subtile_8__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_8__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_8__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_8__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_8__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_8__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_8__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_9__pin_f2a_i_0_(cbx_2__7__4_top_grid_bottom_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_9__pin_sc_in_0_(grid_io_top_8__8__undriven_bottom_width_0_height_0_subtile_9__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_9__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_9__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_9__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_9__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_9__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_9__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_10__pin_f2a_i_0_(cbx_2__7__4_top_grid_bottom_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_10__pin_sc_in_0_(grid_io_top_8__8__undriven_bottom_width_0_height_0_subtile_10__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_10__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_10__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_10__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_10__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_10__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_10__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_11__pin_f2a_i_0_(cbx_2__7__4_top_grid_bottom_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_11__pin_sc_in_0_(grid_io_top_8__8__undriven_bottom_width_0_height_0_subtile_11__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_11__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_11__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_11__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_11__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_11__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_11__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_12__pin_f2a_i_0_(cbx_2__7__4_top_grid_bottom_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_12__pin_sc_in_0_(grid_io_top_8__8__undriven_bottom_width_0_height_0_subtile_12__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_12__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_12__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_12__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_12__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_12__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_12__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_13__pin_f2a_i_0_(cbx_2__7__4_top_grid_bottom_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_13__pin_sc_in_0_(grid_io_top_8__8__undriven_bottom_width_0_height_0_subtile_13__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_13__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_13__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_13__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_13__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_13__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_13__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_14__pin_f2a_i_0_(cbx_2__7__4_top_grid_bottom_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_14__pin_sc_in_0_(grid_io_top_8__8__undriven_bottom_width_0_height_0_subtile_14__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_14__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_14__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_14__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_14__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_14__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_14__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_15__pin_f2a_i_0_(cbx_2__7__4_top_grid_bottom_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_15__pin_sc_in_0_(grid_io_top_8__8__undriven_bottom_width_0_height_0_subtile_15__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_15__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_15__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_15__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_15__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_15__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_15__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_16__pin_f2a_i_0_(cbx_2__7__4_top_grid_bottom_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_16__pin_sc_in_0_(grid_io_top_8__8__undriven_bottom_width_0_height_0_subtile_16__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_16__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_16__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_16__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_16__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_16__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_16__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_17__pin_f2a_i_0_(cbx_2__7__4_top_grid_bottom_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_17__pin_sc_in_0_(grid_io_top_8__8__undriven_bottom_width_0_height_0_subtile_17__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_17__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_17__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_17__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_17__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_17__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_17__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_18__pin_f2a_i_0_(cbx_2__7__4_top_grid_bottom_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_18__pin_sc_in_0_(grid_io_top_8__8__undriven_bottom_width_0_height_0_subtile_18__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_18__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_18__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_18__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_18__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_18__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_18__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_19__pin_f2a_i_0_(cbx_2__7__4_top_grid_bottom_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_19__pin_sc_in_0_(grid_io_top_8__8__undriven_bottom_width_0_height_0_subtile_19__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_19__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_19__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_19__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_19__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_19__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_19__pin_clk_3_(clk[3]),
		.ccff_head(cbx_2__7__4_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_io_top_8__8__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_1__pin_sc_out_0_(grid_io_top_8__8__undriven_bottom_width_0_height_0_subtile_1__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_2__pin_sc_out_0_(grid_io_top_8__8__undriven_bottom_width_0_height_0_subtile_2__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_3__pin_sc_out_0_(grid_io_top_8__8__undriven_bottom_width_0_height_0_subtile_3__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_4__pin_sc_out_0_(grid_io_top_8__8__undriven_bottom_width_0_height_0_subtile_4__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_5__pin_sc_out_0_(grid_io_top_8__8__undriven_bottom_width_0_height_0_subtile_5__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_6__pin_sc_out_0_(grid_io_top_8__8__undriven_bottom_width_0_height_0_subtile_6__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_7__pin_sc_out_0_(grid_io_top_8__8__undriven_bottom_width_0_height_0_subtile_7__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_8__pin_sc_out_0_(grid_io_top_8__8__undriven_bottom_width_0_height_0_subtile_8__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_9__pin_sc_out_0_(grid_io_top_8__8__undriven_bottom_width_0_height_0_subtile_9__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_10__pin_sc_out_0_(grid_io_top_8__8__undriven_bottom_width_0_height_0_subtile_10__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_11__pin_sc_out_0_(grid_io_top_8__8__undriven_bottom_width_0_height_0_subtile_11__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_12__pin_sc_out_0_(grid_io_top_8__8__undriven_bottom_width_0_height_0_subtile_12__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_13__pin_sc_out_0_(grid_io_top_8__8__undriven_bottom_width_0_height_0_subtile_13__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_14__pin_sc_out_0_(grid_io_top_8__8__undriven_bottom_width_0_height_0_subtile_14__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_15__pin_sc_out_0_(grid_io_top_8__8__undriven_bottom_width_0_height_0_subtile_15__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_16__pin_sc_out_0_(grid_io_top_8__8__undriven_bottom_width_0_height_0_subtile_16__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_17__pin_sc_out_0_(grid_io_top_8__8__undriven_bottom_width_0_height_0_subtile_17__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_18__pin_sc_out_0_(grid_io_top_8__8__undriven_bottom_width_0_height_0_subtile_18__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_19__pin_sc_out_0_(grid_io_top_8__8__undriven_bottom_width_0_height_0_subtile_19__pin_sc_out_0_),
		.ccff_tail(grid_io_top_6_ccff_tail));

	grid_io_top grid_io_top_9__8_ (
		.test_en(test_en),
		.scan_mode(scan_mode),
		.scan_clk(scan_clk),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.CFG_DONE(CFG_DONE),
		.gfpga_pad_QL_PREIO_A2F(gfpga_pad_QL_PREIO_A2F[300:319]),
		.gfpga_pad_QL_PREIO_F2A(gfpga_pad_QL_PREIO_F2A[300:319]),
		.gfpga_pad_QL_PREIO_F2A_DEF0(gfpga_pad_QL_PREIO_F2A_DEF0[300:319]),
		.gfpga_pad_QL_PREIO_F2A_DEF1(gfpga_pad_QL_PREIO_F2A_DEF1[300:319]),
		.gfpga_pad_QL_PREIO_F2A_CLK(gfpga_pad_QL_PREIO_F2A_CLK[300:319]),
		.bottom_width_0_height_0_subtile_0__pin_f2a_i_0_(cbx_2__7__5_top_grid_bottom_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_in_0_(grid_io_top_9__8__undriven_bottom_width_0_height_0_subtile_0__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_1__pin_f2a_i_0_(cbx_2__7__5_top_grid_bottom_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_1__pin_sc_in_0_(grid_io_top_9__8__undriven_bottom_width_0_height_0_subtile_1__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_1__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_1__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_1__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_1__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_1__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_1__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_2__pin_f2a_i_0_(cbx_2__7__5_top_grid_bottom_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_2__pin_sc_in_0_(grid_io_top_9__8__undriven_bottom_width_0_height_0_subtile_2__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_2__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_2__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_2__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_2__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_2__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_2__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_3__pin_f2a_i_0_(cbx_2__7__5_top_grid_bottom_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_3__pin_sc_in_0_(grid_io_top_9__8__undriven_bottom_width_0_height_0_subtile_3__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_3__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_3__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_3__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_3__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_3__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_3__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_4__pin_f2a_i_0_(cbx_2__7__5_top_grid_bottom_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_4__pin_sc_in_0_(grid_io_top_9__8__undriven_bottom_width_0_height_0_subtile_4__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_4__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_4__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_4__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_4__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_4__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_4__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_5__pin_f2a_i_0_(cbx_2__7__5_top_grid_bottom_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_5__pin_sc_in_0_(grid_io_top_9__8__undriven_bottom_width_0_height_0_subtile_5__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_5__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_5__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_5__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_5__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_5__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_5__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_6__pin_f2a_i_0_(cbx_2__7__5_top_grid_bottom_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_6__pin_sc_in_0_(grid_io_top_9__8__undriven_bottom_width_0_height_0_subtile_6__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_6__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_6__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_6__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_6__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_6__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_6__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_7__pin_f2a_i_0_(cbx_2__7__5_top_grid_bottom_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_7__pin_sc_in_0_(grid_io_top_9__8__undriven_bottom_width_0_height_0_subtile_7__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_7__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_7__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_7__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_7__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_7__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_7__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_8__pin_f2a_i_0_(cbx_2__7__5_top_grid_bottom_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_8__pin_sc_in_0_(grid_io_top_9__8__undriven_bottom_width_0_height_0_subtile_8__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_8__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_8__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_8__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_8__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_8__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_8__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_9__pin_f2a_i_0_(cbx_2__7__5_top_grid_bottom_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_9__pin_sc_in_0_(grid_io_top_9__8__undriven_bottom_width_0_height_0_subtile_9__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_9__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_9__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_9__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_9__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_9__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_9__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_10__pin_f2a_i_0_(cbx_2__7__5_top_grid_bottom_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_10__pin_sc_in_0_(grid_io_top_9__8__undriven_bottom_width_0_height_0_subtile_10__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_10__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_10__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_10__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_10__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_10__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_10__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_11__pin_f2a_i_0_(cbx_2__7__5_top_grid_bottom_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_11__pin_sc_in_0_(grid_io_top_9__8__undriven_bottom_width_0_height_0_subtile_11__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_11__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_11__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_11__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_11__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_11__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_11__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_12__pin_f2a_i_0_(cbx_2__7__5_top_grid_bottom_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_12__pin_sc_in_0_(grid_io_top_9__8__undriven_bottom_width_0_height_0_subtile_12__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_12__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_12__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_12__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_12__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_12__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_12__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_13__pin_f2a_i_0_(cbx_2__7__5_top_grid_bottom_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_13__pin_sc_in_0_(grid_io_top_9__8__undriven_bottom_width_0_height_0_subtile_13__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_13__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_13__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_13__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_13__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_13__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_13__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_14__pin_f2a_i_0_(cbx_2__7__5_top_grid_bottom_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_14__pin_sc_in_0_(grid_io_top_9__8__undriven_bottom_width_0_height_0_subtile_14__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_14__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_14__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_14__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_14__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_14__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_14__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_15__pin_f2a_i_0_(cbx_2__7__5_top_grid_bottom_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_15__pin_sc_in_0_(grid_io_top_9__8__undriven_bottom_width_0_height_0_subtile_15__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_15__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_15__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_15__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_15__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_15__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_15__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_16__pin_f2a_i_0_(cbx_2__7__5_top_grid_bottom_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_16__pin_sc_in_0_(grid_io_top_9__8__undriven_bottom_width_0_height_0_subtile_16__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_16__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_16__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_16__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_16__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_16__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_16__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_17__pin_f2a_i_0_(cbx_2__7__5_top_grid_bottom_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_17__pin_sc_in_0_(grid_io_top_9__8__undriven_bottom_width_0_height_0_subtile_17__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_17__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_17__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_17__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_17__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_17__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_17__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_18__pin_f2a_i_0_(cbx_2__7__5_top_grid_bottom_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_18__pin_sc_in_0_(grid_io_top_9__8__undriven_bottom_width_0_height_0_subtile_18__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_18__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_18__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_18__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_18__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_18__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_18__pin_clk_3_(clk[3]),
		.bottom_width_0_height_0_subtile_19__pin_f2a_i_0_(cbx_2__7__5_top_grid_bottom_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.bottom_width_0_height_0_subtile_19__pin_sc_in_0_(grid_io_top_9__8__undriven_bottom_width_0_height_0_subtile_19__pin_sc_in_0_),
		.bottom_width_0_height_0_subtile_19__pin_global_reset_0_(global_reset),
		.bottom_width_0_height_0_subtile_19__pin_scan_reset_0_(scan_reset),
		.bottom_width_0_height_0_subtile_19__pin_clk_0_(clk[0]),
		.bottom_width_0_height_0_subtile_19__pin_clk_1_(clk[1]),
		.bottom_width_0_height_0_subtile_19__pin_clk_2_(clk[2]),
		.bottom_width_0_height_0_subtile_19__pin_clk_3_(clk[3]),
		.ccff_head(cby_9__1__1_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_io_top_9__8__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_1__pin_sc_out_0_(grid_io_top_9__8__undriven_bottom_width_0_height_0_subtile_1__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_2__pin_sc_out_0_(grid_io_top_9__8__undriven_bottom_width_0_height_0_subtile_2__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_3__pin_sc_out_0_(grid_io_top_9__8__undriven_bottom_width_0_height_0_subtile_3__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_4__pin_sc_out_0_(grid_io_top_9__8__undriven_bottom_width_0_height_0_subtile_4__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_5__pin_sc_out_0_(grid_io_top_9__8__undriven_bottom_width_0_height_0_subtile_5__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_6__pin_sc_out_0_(grid_io_top_9__8__undriven_bottom_width_0_height_0_subtile_6__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_7__pin_sc_out_0_(grid_io_top_9__8__undriven_bottom_width_0_height_0_subtile_7__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_8__pin_sc_out_0_(grid_io_top_9__8__undriven_bottom_width_0_height_0_subtile_8__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_9__pin_sc_out_0_(grid_io_top_9__8__undriven_bottom_width_0_height_0_subtile_9__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_10__pin_sc_out_0_(grid_io_top_9__8__undriven_bottom_width_0_height_0_subtile_10__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_11__pin_sc_out_0_(grid_io_top_9__8__undriven_bottom_width_0_height_0_subtile_11__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_12__pin_sc_out_0_(grid_io_top_9__8__undriven_bottom_width_0_height_0_subtile_12__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_13__pin_sc_out_0_(grid_io_top_9__8__undriven_bottom_width_0_height_0_subtile_13__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_14__pin_sc_out_0_(grid_io_top_9__8__undriven_bottom_width_0_height_0_subtile_14__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_15__pin_sc_out_0_(grid_io_top_9__8__undriven_bottom_width_0_height_0_subtile_15__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_16__pin_sc_out_0_(grid_io_top_9__8__undriven_bottom_width_0_height_0_subtile_16__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_17__pin_sc_out_0_(grid_io_top_9__8__undriven_bottom_width_0_height_0_subtile_17__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_18__pin_sc_out_0_(grid_io_top_9__8__undriven_bottom_width_0_height_0_subtile_18__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.bottom_width_0_height_0_subtile_19__pin_sc_out_0_(grid_io_top_9__8__undriven_bottom_width_0_height_0_subtile_19__pin_sc_out_0_),
		.ccff_tail(grid_io_top_7_ccff_tail));

	grid_dsp grid_dsp_4__2_ (
		.test_en(test_en),
		.scan_mode(scan_mode),
		.scan_clk(scan_clk),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_dsp_4__2__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_1_(grid_dsp_4__2__undriven_top_width_0_height_0_subtile_0__pin_sc_in_1_),
		.top_width_0_height_0_subtile_0__pin_sc_in_2_(grid_dsp_4__2__undriven_top_width_0_height_0_subtile_0__pin_sc_in_2_),
		.top_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_0__pin_a_i_2_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_a_i_2_),
		.right_width_0_height_0_subtile_0__pin_a_i_3_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_a_i_3_),
		.right_width_0_height_0_subtile_0__pin_a_i_4_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_a_i_4_),
		.right_width_0_height_0_subtile_0__pin_a_i_5_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_a_i_5_),
		.right_width_0_height_0_subtile_0__pin_a_i_6_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_a_i_6_),
		.right_width_0_height_0_subtile_0__pin_a_i_7_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_a_i_7_),
		.right_width_0_height_0_subtile_0__pin_acc_fir_i_1_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_acc_fir_i_1_),
		.right_width_0_height_0_subtile_0__pin_acc_fir_i_2_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_acc_fir_i_2_),
		.right_width_0_height_0_subtile_0__pin_b_i_0_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_b_i_0_),
		.right_width_0_height_0_subtile_0__pin_b_i_1_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_b_i_1_),
		.right_width_0_height_0_subtile_0__pin_b_i_2_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_b_i_2_),
		.right_width_0_height_0_subtile_0__pin_b_i_3_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_b_i_3_),
		.right_width_0_height_0_subtile_0__pin_b_i_4_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_b_i_4_),
		.right_width_0_height_0_subtile_0__pin_b_i_5_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_b_i_5_),
		.right_width_0_height_0_subtile_0__pin_unsigned_a_0_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_unsigned_a_0_),
		.right_width_0_height_0_subtile_0__pin_round_0_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_round_0_),
		.right_width_0_height_1_subtile_0__pin_a_i_8_(cby_4__3__0_left_grid_right_width_0_height_1_subtile_0__pin_a_i_8_),
		.right_width_0_height_1_subtile_0__pin_a_i_9_(cby_4__3__0_left_grid_right_width_0_height_1_subtile_0__pin_a_i_9_),
		.right_width_0_height_1_subtile_0__pin_a_i_10_(cby_4__3__0_left_grid_right_width_0_height_1_subtile_0__pin_a_i_10_),
		.right_width_0_height_1_subtile_0__pin_a_i_11_(cby_4__3__0_left_grid_right_width_0_height_1_subtile_0__pin_a_i_11_),
		.right_width_0_height_1_subtile_0__pin_a_i_12_(cby_4__3__0_left_grid_right_width_0_height_1_subtile_0__pin_a_i_12_),
		.right_width_0_height_1_subtile_0__pin_a_i_13_(cby_4__3__0_left_grid_right_width_0_height_1_subtile_0__pin_a_i_13_),
		.right_width_0_height_1_subtile_0__pin_acc_fir_i_3_(cby_4__3__0_left_grid_right_width_0_height_1_subtile_0__pin_acc_fir_i_3_),
		.right_width_0_height_1_subtile_0__pin_acc_fir_i_4_(cby_4__3__0_left_grid_right_width_0_height_1_subtile_0__pin_acc_fir_i_4_),
		.right_width_0_height_1_subtile_0__pin_b_i_6_(cby_4__3__0_left_grid_right_width_0_height_1_subtile_0__pin_b_i_6_),
		.right_width_0_height_1_subtile_0__pin_b_i_7_(cby_4__3__0_left_grid_right_width_0_height_1_subtile_0__pin_b_i_7_),
		.right_width_0_height_1_subtile_0__pin_b_i_8_(cby_4__3__0_left_grid_right_width_0_height_1_subtile_0__pin_b_i_8_),
		.right_width_0_height_1_subtile_0__pin_b_i_9_(cby_4__3__0_left_grid_right_width_0_height_1_subtile_0__pin_b_i_9_),
		.right_width_0_height_1_subtile_0__pin_b_i_10_(cby_4__3__0_left_grid_right_width_0_height_1_subtile_0__pin_b_i_10_),
		.right_width_0_height_1_subtile_0__pin_b_i_11_(cby_4__3__0_left_grid_right_width_0_height_1_subtile_0__pin_b_i_11_),
		.right_width_0_height_1_subtile_0__pin_unsigned_b_0_(cby_4__3__0_left_grid_right_width_0_height_1_subtile_0__pin_unsigned_b_0_),
		.right_width_0_height_1_subtile_0__pin_subtract_0_(cby_4__3__0_left_grid_right_width_0_height_1_subtile_0__pin_subtract_0_),
		.right_width_0_height_2_subtile_0__pin_a_i_14_(cby_4__4__0_left_grid_right_width_0_height_2_subtile_0__pin_a_i_14_),
		.right_width_0_height_2_subtile_0__pin_a_i_15_(cby_4__4__0_left_grid_right_width_0_height_2_subtile_0__pin_a_i_15_),
		.right_width_0_height_2_subtile_0__pin_a_i_16_(cby_4__4__0_left_grid_right_width_0_height_2_subtile_0__pin_a_i_16_),
		.right_width_0_height_2_subtile_0__pin_a_i_17_(cby_4__4__0_left_grid_right_width_0_height_2_subtile_0__pin_a_i_17_),
		.right_width_0_height_2_subtile_0__pin_a_i_18_(cby_4__4__0_left_grid_right_width_0_height_2_subtile_0__pin_a_i_18_),
		.right_width_0_height_2_subtile_0__pin_a_i_19_(cby_4__4__0_left_grid_right_width_0_height_2_subtile_0__pin_a_i_19_),
		.right_width_0_height_2_subtile_0__pin_acc_fir_i_5_(cby_4__4__0_left_grid_right_width_0_height_2_subtile_0__pin_acc_fir_i_5_),
		.right_width_0_height_2_subtile_0__pin_b_i_12_(cby_4__4__0_left_grid_right_width_0_height_2_subtile_0__pin_b_i_12_),
		.right_width_0_height_2_subtile_0__pin_b_i_13_(cby_4__4__0_left_grid_right_width_0_height_2_subtile_0__pin_b_i_13_),
		.right_width_0_height_2_subtile_0__pin_b_i_14_(cby_4__4__0_left_grid_right_width_0_height_2_subtile_0__pin_b_i_14_),
		.right_width_0_height_2_subtile_0__pin_b_i_15_(cby_4__4__0_left_grid_right_width_0_height_2_subtile_0__pin_b_i_15_),
		.right_width_0_height_2_subtile_0__pin_b_i_16_(cby_4__4__0_left_grid_right_width_0_height_2_subtile_0__pin_b_i_16_),
		.right_width_0_height_2_subtile_0__pin_b_i_17_(cby_4__4__0_left_grid_right_width_0_height_2_subtile_0__pin_b_i_17_),
		.right_width_0_height_2_subtile_0__pin_load_acc_0_(cby_4__4__0_left_grid_right_width_0_height_2_subtile_0__pin_load_acc_0_),
		.right_width_0_height_2_subtile_0__pin_saturate_enable_0_(cby_4__4__0_left_grid_right_width_0_height_2_subtile_0__pin_saturate_enable_0_),
		.bottom_width_0_height_0_subtile_0__pin_a_i_0_(cbx_4__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_a_i_0_),
		.bottom_width_0_height_0_subtile_0__pin_a_i_1_(cbx_4__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_a_i_1_),
		.bottom_width_0_height_0_subtile_0__pin_acc_fir_i_0_(cbx_4__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_acc_fir_i_0_),
		.bottom_width_0_height_0_subtile_0__pin_lreset_0_(cbx_4__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_lreset_0_),
		.bottom_width_0_height_0_subtile_0__pin_feedback_0_(cbx_4__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_feedback_0_),
		.bottom_width_0_height_0_subtile_0__pin_feedback_1_(cbx_4__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_feedback_1_),
		.bottom_width_0_height_0_subtile_0__pin_feedback_2_(cbx_4__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_feedback_2_),
		.bottom_width_0_height_0_subtile_0__pin_shift_right_0_(cbx_4__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_shift_right_0_),
		.bottom_width_0_height_0_subtile_0__pin_shift_right_1_(cbx_4__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_shift_right_1_),
		.bottom_width_0_height_0_subtile_0__pin_shift_right_2_(cbx_4__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_shift_right_2_),
		.bottom_width_0_height_0_subtile_0__pin_shift_right_3_(cbx_4__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_shift_right_3_),
		.bottom_width_0_height_0_subtile_0__pin_shift_right_4_(cbx_4__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_shift_right_4_),
		.bottom_width_0_height_0_subtile_0__pin_shift_right_5_(cbx_4__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_shift_right_5_),
		.ccff_head(cby_4__2__0_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_z_o_7_(grid_dsp_0_right_width_0_height_0_subtile_0__pin_z_o_7_),
		.right_width_0_height_0_subtile_0__pin_z_o_8_(grid_dsp_0_right_width_0_height_0_subtile_0__pin_z_o_8_),
		.right_width_0_height_0_subtile_0__pin_z_o_9_(grid_dsp_0_right_width_0_height_0_subtile_0__pin_z_o_9_),
		.right_width_0_height_0_subtile_0__pin_z_o_10_(grid_dsp_0_right_width_0_height_0_subtile_0__pin_z_o_10_),
		.right_width_0_height_0_subtile_0__pin_z_o_11_(grid_dsp_0_right_width_0_height_0_subtile_0__pin_z_o_11_),
		.right_width_0_height_0_subtile_0__pin_z_o_12_(grid_dsp_0_right_width_0_height_0_subtile_0__pin_z_o_12_),
		.right_width_0_height_0_subtile_0__pin_z_o_13_(grid_dsp_0_right_width_0_height_0_subtile_0__pin_z_o_13_),
		.right_width_0_height_0_subtile_0__pin_z_o_14_(grid_dsp_0_right_width_0_height_0_subtile_0__pin_z_o_14_),
		.right_width_0_height_0_subtile_0__pin_z_o_15_(grid_dsp_0_right_width_0_height_0_subtile_0__pin_z_o_15_),
		.right_width_0_height_0_subtile_0__pin_dly_b_o_0_(grid_dsp_0_right_width_0_height_0_subtile_0__pin_dly_b_o_0_),
		.right_width_0_height_0_subtile_0__pin_dly_b_o_1_(grid_dsp_0_right_width_0_height_0_subtile_0__pin_dly_b_o_1_),
		.right_width_0_height_0_subtile_0__pin_dly_b_o_2_(grid_dsp_0_right_width_0_height_0_subtile_0__pin_dly_b_o_2_),
		.right_width_0_height_0_subtile_0__pin_dly_b_o_3_(grid_dsp_0_right_width_0_height_0_subtile_0__pin_dly_b_o_3_),
		.right_width_0_height_0_subtile_0__pin_dly_b_o_4_(grid_dsp_0_right_width_0_height_0_subtile_0__pin_dly_b_o_4_),
		.right_width_0_height_0_subtile_0__pin_dly_b_o_5_(grid_dsp_0_right_width_0_height_0_subtile_0__pin_dly_b_o_5_),
		.right_width_0_height_1_subtile_0__pin_z_o_16_(grid_dsp_0_right_width_0_height_1_subtile_0__pin_z_o_16_),
		.right_width_0_height_1_subtile_0__pin_z_o_17_(grid_dsp_0_right_width_0_height_1_subtile_0__pin_z_o_17_),
		.right_width_0_height_1_subtile_0__pin_z_o_18_(grid_dsp_0_right_width_0_height_1_subtile_0__pin_z_o_18_),
		.right_width_0_height_1_subtile_0__pin_z_o_19_(grid_dsp_0_right_width_0_height_1_subtile_0__pin_z_o_19_),
		.right_width_0_height_1_subtile_0__pin_z_o_20_(grid_dsp_0_right_width_0_height_1_subtile_0__pin_z_o_20_),
		.right_width_0_height_1_subtile_0__pin_z_o_21_(grid_dsp_0_right_width_0_height_1_subtile_0__pin_z_o_21_),
		.right_width_0_height_1_subtile_0__pin_z_o_22_(grid_dsp_0_right_width_0_height_1_subtile_0__pin_z_o_22_),
		.right_width_0_height_1_subtile_0__pin_z_o_23_(grid_dsp_0_right_width_0_height_1_subtile_0__pin_z_o_23_),
		.right_width_0_height_1_subtile_0__pin_z_o_24_(grid_dsp_0_right_width_0_height_1_subtile_0__pin_z_o_24_),
		.right_width_0_height_1_subtile_0__pin_z_o_25_(grid_dsp_0_right_width_0_height_1_subtile_0__pin_z_o_25_),
		.right_width_0_height_1_subtile_0__pin_z_o_26_(grid_dsp_0_right_width_0_height_1_subtile_0__pin_z_o_26_),
		.right_width_0_height_1_subtile_0__pin_dly_b_o_6_(grid_dsp_0_right_width_0_height_1_subtile_0__pin_dly_b_o_6_),
		.right_width_0_height_1_subtile_0__pin_dly_b_o_7_(grid_dsp_0_right_width_0_height_1_subtile_0__pin_dly_b_o_7_),
		.right_width_0_height_1_subtile_0__pin_dly_b_o_8_(grid_dsp_0_right_width_0_height_1_subtile_0__pin_dly_b_o_8_),
		.right_width_0_height_1_subtile_0__pin_dly_b_o_9_(grid_dsp_0_right_width_0_height_1_subtile_0__pin_dly_b_o_9_),
		.right_width_0_height_1_subtile_0__pin_dly_b_o_10_(grid_dsp_0_right_width_0_height_1_subtile_0__pin_dly_b_o_10_),
		.right_width_0_height_1_subtile_0__pin_dly_b_o_11_(grid_dsp_0_right_width_0_height_1_subtile_0__pin_dly_b_o_11_),
		.right_width_0_height_2_subtile_0__pin_z_o_27_(grid_dsp_0_right_width_0_height_2_subtile_0__pin_z_o_27_),
		.right_width_0_height_2_subtile_0__pin_z_o_28_(grid_dsp_0_right_width_0_height_2_subtile_0__pin_z_o_28_),
		.right_width_0_height_2_subtile_0__pin_z_o_29_(grid_dsp_0_right_width_0_height_2_subtile_0__pin_z_o_29_),
		.right_width_0_height_2_subtile_0__pin_z_o_30_(grid_dsp_0_right_width_0_height_2_subtile_0__pin_z_o_30_),
		.right_width_0_height_2_subtile_0__pin_z_o_31_(grid_dsp_0_right_width_0_height_2_subtile_0__pin_z_o_31_),
		.right_width_0_height_2_subtile_0__pin_z_o_32_(grid_dsp_0_right_width_0_height_2_subtile_0__pin_z_o_32_),
		.right_width_0_height_2_subtile_0__pin_z_o_33_(grid_dsp_0_right_width_0_height_2_subtile_0__pin_z_o_33_),
		.right_width_0_height_2_subtile_0__pin_z_o_34_(grid_dsp_0_right_width_0_height_2_subtile_0__pin_z_o_34_),
		.right_width_0_height_2_subtile_0__pin_z_o_35_(grid_dsp_0_right_width_0_height_2_subtile_0__pin_z_o_35_),
		.right_width_0_height_2_subtile_0__pin_z_o_36_(grid_dsp_0_right_width_0_height_2_subtile_0__pin_z_o_36_),
		.right_width_0_height_2_subtile_0__pin_z_o_37_(grid_dsp_0_right_width_0_height_2_subtile_0__pin_z_o_37_),
		.right_width_0_height_2_subtile_0__pin_dly_b_o_12_(grid_dsp_0_right_width_0_height_2_subtile_0__pin_dly_b_o_12_),
		.right_width_0_height_2_subtile_0__pin_dly_b_o_13_(grid_dsp_0_right_width_0_height_2_subtile_0__pin_dly_b_o_13_),
		.right_width_0_height_2_subtile_0__pin_dly_b_o_14_(grid_dsp_0_right_width_0_height_2_subtile_0__pin_dly_b_o_14_),
		.right_width_0_height_2_subtile_0__pin_dly_b_o_15_(grid_dsp_0_right_width_0_height_2_subtile_0__pin_dly_b_o_15_),
		.right_width_0_height_2_subtile_0__pin_dly_b_o_16_(grid_dsp_0_right_width_0_height_2_subtile_0__pin_dly_b_o_16_),
		.right_width_0_height_2_subtile_0__pin_dly_b_o_17_(grid_dsp_0_right_width_0_height_2_subtile_0__pin_dly_b_o_17_),
		.bottom_width_0_height_0_subtile_0__pin_z_o_0_(grid_dsp_0_bottom_width_0_height_0_subtile_0__pin_z_o_0_),
		.bottom_width_0_height_0_subtile_0__pin_z_o_1_(grid_dsp_0_bottom_width_0_height_0_subtile_0__pin_z_o_1_),
		.bottom_width_0_height_0_subtile_0__pin_z_o_2_(grid_dsp_0_bottom_width_0_height_0_subtile_0__pin_z_o_2_),
		.bottom_width_0_height_0_subtile_0__pin_z_o_3_(grid_dsp_0_bottom_width_0_height_0_subtile_0__pin_z_o_3_),
		.bottom_width_0_height_0_subtile_0__pin_z_o_4_(grid_dsp_0_bottom_width_0_height_0_subtile_0__pin_z_o_4_),
		.bottom_width_0_height_0_subtile_0__pin_z_o_5_(grid_dsp_0_bottom_width_0_height_0_subtile_0__pin_z_o_5_),
		.bottom_width_0_height_0_subtile_0__pin_z_o_6_(grid_dsp_0_bottom_width_0_height_0_subtile_0__pin_z_o_6_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_dsp_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_1_(grid_dsp_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_1_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_2_(grid_dsp_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_2_),
		.ccff_tail(grid_dsp_0_ccff_tail));

	grid_dsp grid_dsp_4__5_ (
		.test_en(test_en),
		.scan_mode(scan_mode),
		.scan_clk(scan_clk),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_dsp_4__5__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_1_(grid_dsp_4__5__undriven_top_width_0_height_0_subtile_0__pin_sc_in_1_),
		.top_width_0_height_0_subtile_0__pin_sc_in_2_(grid_dsp_4__5__undriven_top_width_0_height_0_subtile_0__pin_sc_in_2_),
		.top_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.top_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.top_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.top_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.top_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.top_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.right_width_0_height_0_subtile_0__pin_a_i_2_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_a_i_2_),
		.right_width_0_height_0_subtile_0__pin_a_i_3_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_a_i_3_),
		.right_width_0_height_0_subtile_0__pin_a_i_4_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_a_i_4_),
		.right_width_0_height_0_subtile_0__pin_a_i_5_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_a_i_5_),
		.right_width_0_height_0_subtile_0__pin_a_i_6_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_a_i_6_),
		.right_width_0_height_0_subtile_0__pin_a_i_7_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_a_i_7_),
		.right_width_0_height_0_subtile_0__pin_acc_fir_i_1_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_acc_fir_i_1_),
		.right_width_0_height_0_subtile_0__pin_acc_fir_i_2_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_acc_fir_i_2_),
		.right_width_0_height_0_subtile_0__pin_b_i_0_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_b_i_0_),
		.right_width_0_height_0_subtile_0__pin_b_i_1_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_b_i_1_),
		.right_width_0_height_0_subtile_0__pin_b_i_2_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_b_i_2_),
		.right_width_0_height_0_subtile_0__pin_b_i_3_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_b_i_3_),
		.right_width_0_height_0_subtile_0__pin_b_i_4_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_b_i_4_),
		.right_width_0_height_0_subtile_0__pin_b_i_5_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_b_i_5_),
		.right_width_0_height_0_subtile_0__pin_unsigned_a_0_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_unsigned_a_0_),
		.right_width_0_height_0_subtile_0__pin_round_0_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_round_0_),
		.right_width_0_height_1_subtile_0__pin_a_i_8_(cby_4__3__1_left_grid_right_width_0_height_1_subtile_0__pin_a_i_8_),
		.right_width_0_height_1_subtile_0__pin_a_i_9_(cby_4__3__1_left_grid_right_width_0_height_1_subtile_0__pin_a_i_9_),
		.right_width_0_height_1_subtile_0__pin_a_i_10_(cby_4__3__1_left_grid_right_width_0_height_1_subtile_0__pin_a_i_10_),
		.right_width_0_height_1_subtile_0__pin_a_i_11_(cby_4__3__1_left_grid_right_width_0_height_1_subtile_0__pin_a_i_11_),
		.right_width_0_height_1_subtile_0__pin_a_i_12_(cby_4__3__1_left_grid_right_width_0_height_1_subtile_0__pin_a_i_12_),
		.right_width_0_height_1_subtile_0__pin_a_i_13_(cby_4__3__1_left_grid_right_width_0_height_1_subtile_0__pin_a_i_13_),
		.right_width_0_height_1_subtile_0__pin_acc_fir_i_3_(cby_4__3__1_left_grid_right_width_0_height_1_subtile_0__pin_acc_fir_i_3_),
		.right_width_0_height_1_subtile_0__pin_acc_fir_i_4_(cby_4__3__1_left_grid_right_width_0_height_1_subtile_0__pin_acc_fir_i_4_),
		.right_width_0_height_1_subtile_0__pin_b_i_6_(cby_4__3__1_left_grid_right_width_0_height_1_subtile_0__pin_b_i_6_),
		.right_width_0_height_1_subtile_0__pin_b_i_7_(cby_4__3__1_left_grid_right_width_0_height_1_subtile_0__pin_b_i_7_),
		.right_width_0_height_1_subtile_0__pin_b_i_8_(cby_4__3__1_left_grid_right_width_0_height_1_subtile_0__pin_b_i_8_),
		.right_width_0_height_1_subtile_0__pin_b_i_9_(cby_4__3__1_left_grid_right_width_0_height_1_subtile_0__pin_b_i_9_),
		.right_width_0_height_1_subtile_0__pin_b_i_10_(cby_4__3__1_left_grid_right_width_0_height_1_subtile_0__pin_b_i_10_),
		.right_width_0_height_1_subtile_0__pin_b_i_11_(cby_4__3__1_left_grid_right_width_0_height_1_subtile_0__pin_b_i_11_),
		.right_width_0_height_1_subtile_0__pin_unsigned_b_0_(cby_4__3__1_left_grid_right_width_0_height_1_subtile_0__pin_unsigned_b_0_),
		.right_width_0_height_1_subtile_0__pin_subtract_0_(cby_4__3__1_left_grid_right_width_0_height_1_subtile_0__pin_subtract_0_),
		.right_width_0_height_2_subtile_0__pin_a_i_14_(cby_4__4__1_left_grid_right_width_0_height_2_subtile_0__pin_a_i_14_),
		.right_width_0_height_2_subtile_0__pin_a_i_15_(cby_4__4__1_left_grid_right_width_0_height_2_subtile_0__pin_a_i_15_),
		.right_width_0_height_2_subtile_0__pin_a_i_16_(cby_4__4__1_left_grid_right_width_0_height_2_subtile_0__pin_a_i_16_),
		.right_width_0_height_2_subtile_0__pin_a_i_17_(cby_4__4__1_left_grid_right_width_0_height_2_subtile_0__pin_a_i_17_),
		.right_width_0_height_2_subtile_0__pin_a_i_18_(cby_4__4__1_left_grid_right_width_0_height_2_subtile_0__pin_a_i_18_),
		.right_width_0_height_2_subtile_0__pin_a_i_19_(cby_4__4__1_left_grid_right_width_0_height_2_subtile_0__pin_a_i_19_),
		.right_width_0_height_2_subtile_0__pin_acc_fir_i_5_(cby_4__4__1_left_grid_right_width_0_height_2_subtile_0__pin_acc_fir_i_5_),
		.right_width_0_height_2_subtile_0__pin_b_i_12_(cby_4__4__1_left_grid_right_width_0_height_2_subtile_0__pin_b_i_12_),
		.right_width_0_height_2_subtile_0__pin_b_i_13_(cby_4__4__1_left_grid_right_width_0_height_2_subtile_0__pin_b_i_13_),
		.right_width_0_height_2_subtile_0__pin_b_i_14_(cby_4__4__1_left_grid_right_width_0_height_2_subtile_0__pin_b_i_14_),
		.right_width_0_height_2_subtile_0__pin_b_i_15_(cby_4__4__1_left_grid_right_width_0_height_2_subtile_0__pin_b_i_15_),
		.right_width_0_height_2_subtile_0__pin_b_i_16_(cby_4__4__1_left_grid_right_width_0_height_2_subtile_0__pin_b_i_16_),
		.right_width_0_height_2_subtile_0__pin_b_i_17_(cby_4__4__1_left_grid_right_width_0_height_2_subtile_0__pin_b_i_17_),
		.right_width_0_height_2_subtile_0__pin_load_acc_0_(cby_4__4__1_left_grid_right_width_0_height_2_subtile_0__pin_load_acc_0_),
		.right_width_0_height_2_subtile_0__pin_saturate_enable_0_(cby_4__4__1_left_grid_right_width_0_height_2_subtile_0__pin_saturate_enable_0_),
		.bottom_width_0_height_0_subtile_0__pin_a_i_0_(cbx_4__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_a_i_0_),
		.bottom_width_0_height_0_subtile_0__pin_a_i_1_(cbx_4__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_a_i_1_),
		.bottom_width_0_height_0_subtile_0__pin_acc_fir_i_0_(cbx_4__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_acc_fir_i_0_),
		.bottom_width_0_height_0_subtile_0__pin_lreset_0_(cbx_4__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_lreset_0_),
		.bottom_width_0_height_0_subtile_0__pin_feedback_0_(cbx_4__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_feedback_0_),
		.bottom_width_0_height_0_subtile_0__pin_feedback_1_(cbx_4__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_feedback_1_),
		.bottom_width_0_height_0_subtile_0__pin_feedback_2_(cbx_4__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_feedback_2_),
		.bottom_width_0_height_0_subtile_0__pin_shift_right_0_(cbx_4__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_shift_right_0_),
		.bottom_width_0_height_0_subtile_0__pin_shift_right_1_(cbx_4__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_shift_right_1_),
		.bottom_width_0_height_0_subtile_0__pin_shift_right_2_(cbx_4__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_shift_right_2_),
		.bottom_width_0_height_0_subtile_0__pin_shift_right_3_(cbx_4__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_shift_right_3_),
		.bottom_width_0_height_0_subtile_0__pin_shift_right_4_(cbx_4__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_shift_right_4_),
		.bottom_width_0_height_0_subtile_0__pin_shift_right_5_(cbx_4__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_shift_right_5_),
		.ccff_head(cby_4__2__1_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_z_o_7_(grid_dsp_1_right_width_0_height_0_subtile_0__pin_z_o_7_),
		.right_width_0_height_0_subtile_0__pin_z_o_8_(grid_dsp_1_right_width_0_height_0_subtile_0__pin_z_o_8_),
		.right_width_0_height_0_subtile_0__pin_z_o_9_(grid_dsp_1_right_width_0_height_0_subtile_0__pin_z_o_9_),
		.right_width_0_height_0_subtile_0__pin_z_o_10_(grid_dsp_1_right_width_0_height_0_subtile_0__pin_z_o_10_),
		.right_width_0_height_0_subtile_0__pin_z_o_11_(grid_dsp_1_right_width_0_height_0_subtile_0__pin_z_o_11_),
		.right_width_0_height_0_subtile_0__pin_z_o_12_(grid_dsp_1_right_width_0_height_0_subtile_0__pin_z_o_12_),
		.right_width_0_height_0_subtile_0__pin_z_o_13_(grid_dsp_1_right_width_0_height_0_subtile_0__pin_z_o_13_),
		.right_width_0_height_0_subtile_0__pin_z_o_14_(grid_dsp_1_right_width_0_height_0_subtile_0__pin_z_o_14_),
		.right_width_0_height_0_subtile_0__pin_z_o_15_(grid_dsp_1_right_width_0_height_0_subtile_0__pin_z_o_15_),
		.right_width_0_height_0_subtile_0__pin_dly_b_o_0_(grid_dsp_1_right_width_0_height_0_subtile_0__pin_dly_b_o_0_),
		.right_width_0_height_0_subtile_0__pin_dly_b_o_1_(grid_dsp_1_right_width_0_height_0_subtile_0__pin_dly_b_o_1_),
		.right_width_0_height_0_subtile_0__pin_dly_b_o_2_(grid_dsp_1_right_width_0_height_0_subtile_0__pin_dly_b_o_2_),
		.right_width_0_height_0_subtile_0__pin_dly_b_o_3_(grid_dsp_1_right_width_0_height_0_subtile_0__pin_dly_b_o_3_),
		.right_width_0_height_0_subtile_0__pin_dly_b_o_4_(grid_dsp_1_right_width_0_height_0_subtile_0__pin_dly_b_o_4_),
		.right_width_0_height_0_subtile_0__pin_dly_b_o_5_(grid_dsp_1_right_width_0_height_0_subtile_0__pin_dly_b_o_5_),
		.right_width_0_height_1_subtile_0__pin_z_o_16_(grid_dsp_1_right_width_0_height_1_subtile_0__pin_z_o_16_),
		.right_width_0_height_1_subtile_0__pin_z_o_17_(grid_dsp_1_right_width_0_height_1_subtile_0__pin_z_o_17_),
		.right_width_0_height_1_subtile_0__pin_z_o_18_(grid_dsp_1_right_width_0_height_1_subtile_0__pin_z_o_18_),
		.right_width_0_height_1_subtile_0__pin_z_o_19_(grid_dsp_1_right_width_0_height_1_subtile_0__pin_z_o_19_),
		.right_width_0_height_1_subtile_0__pin_z_o_20_(grid_dsp_1_right_width_0_height_1_subtile_0__pin_z_o_20_),
		.right_width_0_height_1_subtile_0__pin_z_o_21_(grid_dsp_1_right_width_0_height_1_subtile_0__pin_z_o_21_),
		.right_width_0_height_1_subtile_0__pin_z_o_22_(grid_dsp_1_right_width_0_height_1_subtile_0__pin_z_o_22_),
		.right_width_0_height_1_subtile_0__pin_z_o_23_(grid_dsp_1_right_width_0_height_1_subtile_0__pin_z_o_23_),
		.right_width_0_height_1_subtile_0__pin_z_o_24_(grid_dsp_1_right_width_0_height_1_subtile_0__pin_z_o_24_),
		.right_width_0_height_1_subtile_0__pin_z_o_25_(grid_dsp_1_right_width_0_height_1_subtile_0__pin_z_o_25_),
		.right_width_0_height_1_subtile_0__pin_z_o_26_(grid_dsp_1_right_width_0_height_1_subtile_0__pin_z_o_26_),
		.right_width_0_height_1_subtile_0__pin_dly_b_o_6_(grid_dsp_1_right_width_0_height_1_subtile_0__pin_dly_b_o_6_),
		.right_width_0_height_1_subtile_0__pin_dly_b_o_7_(grid_dsp_1_right_width_0_height_1_subtile_0__pin_dly_b_o_7_),
		.right_width_0_height_1_subtile_0__pin_dly_b_o_8_(grid_dsp_1_right_width_0_height_1_subtile_0__pin_dly_b_o_8_),
		.right_width_0_height_1_subtile_0__pin_dly_b_o_9_(grid_dsp_1_right_width_0_height_1_subtile_0__pin_dly_b_o_9_),
		.right_width_0_height_1_subtile_0__pin_dly_b_o_10_(grid_dsp_1_right_width_0_height_1_subtile_0__pin_dly_b_o_10_),
		.right_width_0_height_1_subtile_0__pin_dly_b_o_11_(grid_dsp_1_right_width_0_height_1_subtile_0__pin_dly_b_o_11_),
		.right_width_0_height_2_subtile_0__pin_z_o_27_(grid_dsp_1_right_width_0_height_2_subtile_0__pin_z_o_27_),
		.right_width_0_height_2_subtile_0__pin_z_o_28_(grid_dsp_1_right_width_0_height_2_subtile_0__pin_z_o_28_),
		.right_width_0_height_2_subtile_0__pin_z_o_29_(grid_dsp_1_right_width_0_height_2_subtile_0__pin_z_o_29_),
		.right_width_0_height_2_subtile_0__pin_z_o_30_(grid_dsp_1_right_width_0_height_2_subtile_0__pin_z_o_30_),
		.right_width_0_height_2_subtile_0__pin_z_o_31_(grid_dsp_1_right_width_0_height_2_subtile_0__pin_z_o_31_),
		.right_width_0_height_2_subtile_0__pin_z_o_32_(grid_dsp_1_right_width_0_height_2_subtile_0__pin_z_o_32_),
		.right_width_0_height_2_subtile_0__pin_z_o_33_(grid_dsp_1_right_width_0_height_2_subtile_0__pin_z_o_33_),
		.right_width_0_height_2_subtile_0__pin_z_o_34_(grid_dsp_1_right_width_0_height_2_subtile_0__pin_z_o_34_),
		.right_width_0_height_2_subtile_0__pin_z_o_35_(grid_dsp_1_right_width_0_height_2_subtile_0__pin_z_o_35_),
		.right_width_0_height_2_subtile_0__pin_z_o_36_(grid_dsp_1_right_width_0_height_2_subtile_0__pin_z_o_36_),
		.right_width_0_height_2_subtile_0__pin_z_o_37_(grid_dsp_1_right_width_0_height_2_subtile_0__pin_z_o_37_),
		.right_width_0_height_2_subtile_0__pin_dly_b_o_12_(grid_dsp_1_right_width_0_height_2_subtile_0__pin_dly_b_o_12_),
		.right_width_0_height_2_subtile_0__pin_dly_b_o_13_(grid_dsp_1_right_width_0_height_2_subtile_0__pin_dly_b_o_13_),
		.right_width_0_height_2_subtile_0__pin_dly_b_o_14_(grid_dsp_1_right_width_0_height_2_subtile_0__pin_dly_b_o_14_),
		.right_width_0_height_2_subtile_0__pin_dly_b_o_15_(grid_dsp_1_right_width_0_height_2_subtile_0__pin_dly_b_o_15_),
		.right_width_0_height_2_subtile_0__pin_dly_b_o_16_(grid_dsp_1_right_width_0_height_2_subtile_0__pin_dly_b_o_16_),
		.right_width_0_height_2_subtile_0__pin_dly_b_o_17_(grid_dsp_1_right_width_0_height_2_subtile_0__pin_dly_b_o_17_),
		.bottom_width_0_height_0_subtile_0__pin_z_o_0_(grid_dsp_1_bottom_width_0_height_0_subtile_0__pin_z_o_0_),
		.bottom_width_0_height_0_subtile_0__pin_z_o_1_(grid_dsp_1_bottom_width_0_height_0_subtile_0__pin_z_o_1_),
		.bottom_width_0_height_0_subtile_0__pin_z_o_2_(grid_dsp_1_bottom_width_0_height_0_subtile_0__pin_z_o_2_),
		.bottom_width_0_height_0_subtile_0__pin_z_o_3_(grid_dsp_1_bottom_width_0_height_0_subtile_0__pin_z_o_3_),
		.bottom_width_0_height_0_subtile_0__pin_z_o_4_(grid_dsp_1_bottom_width_0_height_0_subtile_0__pin_z_o_4_),
		.bottom_width_0_height_0_subtile_0__pin_z_o_5_(grid_dsp_1_bottom_width_0_height_0_subtile_0__pin_z_o_5_),
		.bottom_width_0_height_0_subtile_0__pin_z_o_6_(grid_dsp_1_bottom_width_0_height_0_subtile_0__pin_z_o_6_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_dsp_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_1_(grid_dsp_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_1_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_2_(grid_dsp_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_2_),
		.ccff_tail(grid_dsp_1_ccff_tail));

	grid_bram grid_bram_7__2_ (
		.test_en(test_en),
		.scan_mode(scan_mode),
		.scan_clk(scan_clk),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.top_width_0_height_0_subtile_0__pin_PL_INIT_i_0_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_INIT_i_0_),
		.top_width_0_height_0_subtile_0__pin_PL_ENA_i_0_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_ENA_i_0_),
		.top_width_0_height_0_subtile_0__pin_PL_REN_i_0_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_REN_i_0_),
		.top_width_0_height_0_subtile_0__pin_PL_WEN_i_0_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_WEN_i_0_),
		.top_width_0_height_0_subtile_0__pin_PL_WEN_i_1_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_WEN_i_1_),
		.top_width_0_height_0_subtile_0__pin_PL_ADDR_i_0_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_ADDR_i_0_),
		.top_width_0_height_0_subtile_0__pin_PL_ADDR_i_1_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_ADDR_i_1_),
		.top_width_0_height_0_subtile_0__pin_PL_ADDR_i_2_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_ADDR_i_2_),
		.top_width_0_height_0_subtile_0__pin_PL_ADDR_i_3_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_ADDR_i_3_),
		.top_width_0_height_0_subtile_0__pin_PL_ADDR_i_4_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_ADDR_i_4_),
		.top_width_0_height_0_subtile_0__pin_PL_ADDR_i_5_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_ADDR_i_5_),
		.top_width_0_height_0_subtile_0__pin_PL_ADDR_i_6_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_ADDR_i_6_),
		.top_width_0_height_0_subtile_0__pin_PL_ADDR_i_7_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_ADDR_i_7_),
		.top_width_0_height_0_subtile_0__pin_PL_ADDR_i_8_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_ADDR_i_8_),
		.top_width_0_height_0_subtile_0__pin_PL_ADDR_i_9_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_ADDR_i_9_),
		.top_width_0_height_0_subtile_0__pin_PL_ADDR_i_10_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_ADDR_i_10_),
		.top_width_0_height_0_subtile_0__pin_PL_ADDR_i_11_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_ADDR_i_11_),
		.top_width_0_height_0_subtile_0__pin_PL_ADDR_i_12_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_ADDR_i_12_),
		.top_width_0_height_0_subtile_0__pin_PL_ADDR_i_13_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_ADDR_i_13_),
		.top_width_0_height_0_subtile_0__pin_PL_ADDR_i_14_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_ADDR_i_14_),
		.top_width_0_height_0_subtile_0__pin_PL_ADDR_i_15_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_ADDR_i_15_),
		.top_width_0_height_0_subtile_0__pin_PL_ADDR_i_16_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_ADDR_i_16_),
		.top_width_0_height_0_subtile_0__pin_PL_ADDR_i_17_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_ADDR_i_17_),
		.top_width_0_height_0_subtile_0__pin_PL_ADDR_i_18_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_ADDR_i_18_),
		.top_width_0_height_0_subtile_0__pin_PL_ADDR_i_19_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_ADDR_i_19_),
		.top_width_0_height_0_subtile_0__pin_PL_ADDR_i_20_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_ADDR_i_20_),
		.top_width_0_height_0_subtile_0__pin_PL_ADDR_i_21_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_ADDR_i_21_),
		.top_width_0_height_0_subtile_0__pin_PL_ADDR_i_22_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_ADDR_i_22_),
		.top_width_0_height_0_subtile_0__pin_PL_ADDR_i_23_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_ADDR_i_23_),
		.top_width_0_height_0_subtile_0__pin_PL_ADDR_i_24_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_ADDR_i_24_),
		.top_width_0_height_0_subtile_0__pin_PL_ADDR_i_25_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_ADDR_i_25_),
		.top_width_0_height_0_subtile_0__pin_PL_ADDR_i_26_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_ADDR_i_26_),
		.top_width_0_height_0_subtile_0__pin_PL_ADDR_i_27_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_ADDR_i_27_),
		.top_width_0_height_0_subtile_0__pin_PL_ADDR_i_28_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_ADDR_i_28_),
		.top_width_0_height_0_subtile_0__pin_PL_ADDR_i_29_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_ADDR_i_29_),
		.top_width_0_height_0_subtile_0__pin_PL_ADDR_i_30_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_ADDR_i_30_),
		.top_width_0_height_0_subtile_0__pin_PL_ADDR_i_31_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_ADDR_i_31_),
		.top_width_0_height_0_subtile_0__pin_PL_DATA_i_0_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_DATA_i_0_),
		.top_width_0_height_0_subtile_0__pin_PL_DATA_i_1_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_DATA_i_1_),
		.top_width_0_height_0_subtile_0__pin_PL_DATA_i_2_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_DATA_i_2_),
		.top_width_0_height_0_subtile_0__pin_PL_DATA_i_3_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_DATA_i_3_),
		.top_width_0_height_0_subtile_0__pin_PL_DATA_i_4_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_DATA_i_4_),
		.top_width_0_height_0_subtile_0__pin_PL_DATA_i_5_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_DATA_i_5_),
		.top_width_0_height_0_subtile_0__pin_PL_DATA_i_6_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_DATA_i_6_),
		.top_width_0_height_0_subtile_0__pin_PL_DATA_i_7_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_DATA_i_7_),
		.top_width_0_height_0_subtile_0__pin_PL_DATA_i_8_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_DATA_i_8_),
		.top_width_0_height_0_subtile_0__pin_PL_DATA_i_9_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_DATA_i_9_),
		.top_width_0_height_0_subtile_0__pin_PL_DATA_i_10_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_DATA_i_10_),
		.top_width_0_height_0_subtile_0__pin_PL_DATA_i_11_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_DATA_i_11_),
		.top_width_0_height_0_subtile_0__pin_PL_DATA_i_12_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_DATA_i_12_),
		.top_width_0_height_0_subtile_0__pin_PL_DATA_i_13_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_DATA_i_13_),
		.top_width_0_height_0_subtile_0__pin_PL_DATA_i_14_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_DATA_i_14_),
		.top_width_0_height_0_subtile_0__pin_PL_DATA_i_15_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_DATA_i_15_),
		.top_width_0_height_0_subtile_0__pin_PL_DATA_i_16_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_DATA_i_16_),
		.top_width_0_height_0_subtile_0__pin_PL_DATA_i_17_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_DATA_i_17_),
		.top_width_0_height_0_subtile_0__pin_PL_DATA_i_18_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_DATA_i_18_),
		.top_width_0_height_0_subtile_0__pin_PL_DATA_i_19_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_DATA_i_19_),
		.top_width_0_height_0_subtile_0__pin_PL_DATA_i_20_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_DATA_i_20_),
		.top_width_0_height_0_subtile_0__pin_PL_DATA_i_21_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_DATA_i_21_),
		.top_width_0_height_0_subtile_0__pin_PL_DATA_i_22_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_DATA_i_22_),
		.top_width_0_height_0_subtile_0__pin_PL_DATA_i_23_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_DATA_i_23_),
		.top_width_0_height_0_subtile_0__pin_PL_DATA_i_24_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_DATA_i_24_),
		.top_width_0_height_0_subtile_0__pin_PL_DATA_i_25_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_DATA_i_25_),
		.top_width_0_height_0_subtile_0__pin_PL_DATA_i_26_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_DATA_i_26_),
		.top_width_0_height_0_subtile_0__pin_PL_DATA_i_27_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_DATA_i_27_),
		.top_width_0_height_0_subtile_0__pin_PL_DATA_i_28_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_DATA_i_28_),
		.top_width_0_height_0_subtile_0__pin_PL_DATA_i_29_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_DATA_i_29_),
		.top_width_0_height_0_subtile_0__pin_PL_DATA_i_30_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_DATA_i_30_),
		.top_width_0_height_0_subtile_0__pin_PL_DATA_i_31_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_DATA_i_31_),
		.top_width_0_height_0_subtile_0__pin_PL_DATA_i_32_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_DATA_i_32_),
		.top_width_0_height_0_subtile_0__pin_PL_DATA_i_33_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_DATA_i_33_),
		.top_width_0_height_0_subtile_0__pin_PL_DATA_i_34_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_DATA_i_34_),
		.top_width_0_height_0_subtile_0__pin_PL_DATA_i_35_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_DATA_i_35_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_1_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_sc_in_1_),
		.top_width_0_height_0_subtile_0__pin_sc_in_2_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_sc_in_2_),
		.top_width_0_height_0_subtile_0__pin_sc_in_3_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_sc_in_3_),
		.top_width_0_height_0_subtile_0__pin_sc_in_4_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_sc_in_4_),
		.top_width_0_height_0_subtile_0__pin_sc_in_5_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_sc_in_5_),
		.top_width_0_height_0_subtile_0__pin_PL_CLK_i_0_(grid_bram_7__2__undriven_top_width_0_height_0_subtile_0__pin_PL_CLK_i_0_),
		.right_width_0_height_0_subtile_0__pin_ADDR_A1_i_2_(cby_7__2__0_left_grid_right_width_0_height_0_subtile_0__pin_ADDR_A1_i_2_),
		.right_width_0_height_0_subtile_0__pin_ADDR_A1_i_3_(cby_7__2__0_left_grid_right_width_0_height_0_subtile_0__pin_ADDR_A1_i_3_),
		.right_width_0_height_0_subtile_0__pin_ADDR_A1_i_4_(cby_7__2__0_left_grid_right_width_0_height_0_subtile_0__pin_ADDR_A1_i_4_),
		.right_width_0_height_0_subtile_0__pin_ADDR_A1_i_5_(cby_7__2__0_left_grid_right_width_0_height_0_subtile_0__pin_ADDR_A1_i_5_),
		.right_width_0_height_0_subtile_0__pin_WDATA_B1_i_1_(cby_7__2__0_left_grid_right_width_0_height_0_subtile_0__pin_WDATA_B1_i_1_),
		.right_width_0_height_0_subtile_0__pin_WDATA_B1_i_2_(cby_7__2__0_left_grid_right_width_0_height_0_subtile_0__pin_WDATA_B1_i_2_),
		.right_width_0_height_0_subtile_0__pin_WDATA_B1_i_3_(cby_7__2__0_left_grid_right_width_0_height_0_subtile_0__pin_WDATA_B1_i_3_),
		.right_width_0_height_0_subtile_0__pin_WDATA_B1_i_4_(cby_7__2__0_left_grid_right_width_0_height_0_subtile_0__pin_WDATA_B1_i_4_),
		.right_width_0_height_0_subtile_0__pin_WDATA_B1_i_5_(cby_7__2__0_left_grid_right_width_0_height_0_subtile_0__pin_WDATA_B1_i_5_),
		.right_width_0_height_0_subtile_0__pin_WDATA_B1_i_6_(cby_7__2__0_left_grid_right_width_0_height_0_subtile_0__pin_WDATA_B1_i_6_),
		.right_width_0_height_0_subtile_0__pin_WDATA_B1_i_7_(cby_7__2__0_left_grid_right_width_0_height_0_subtile_0__pin_WDATA_B1_i_7_),
		.right_width_0_height_0_subtile_0__pin_WDATA_B1_i_8_(cby_7__2__0_left_grid_right_width_0_height_0_subtile_0__pin_WDATA_B1_i_8_),
		.right_width_0_height_0_subtile_0__pin_WDATA_B1_i_9_(cby_7__2__0_left_grid_right_width_0_height_0_subtile_0__pin_WDATA_B1_i_9_),
		.right_width_0_height_0_subtile_0__pin_WDATA_B1_i_10_(cby_7__2__0_left_grid_right_width_0_height_0_subtile_0__pin_WDATA_B1_i_10_),
		.right_width_0_height_0_subtile_0__pin_WDATA_B1_i_11_(cby_7__2__0_left_grid_right_width_0_height_0_subtile_0__pin_WDATA_B1_i_11_),
		.right_width_0_height_0_subtile_0__pin_WDATA_B1_i_12_(cby_7__2__0_left_grid_right_width_0_height_0_subtile_0__pin_WDATA_B1_i_12_),
		.right_width_0_height_0_subtile_0__pin_WDATA_B1_i_13_(cby_7__2__0_left_grid_right_width_0_height_0_subtile_0__pin_WDATA_B1_i_13_),
		.right_width_0_height_0_subtile_0__pin_WDATA_B1_i_14_(cby_7__2__0_left_grid_right_width_0_height_0_subtile_0__pin_WDATA_B1_i_14_),
		.right_width_0_height_0_subtile_0__pin_WDATA_B1_i_15_(cby_7__2__0_left_grid_right_width_0_height_0_subtile_0__pin_WDATA_B1_i_15_),
		.right_width_0_height_0_subtile_0__pin_WDATA_B1_i_16_(cby_7__2__0_left_grid_right_width_0_height_0_subtile_0__pin_WDATA_B1_i_16_),
		.right_width_0_height_0_subtile_0__pin_ADDR_B1_i_0_(cby_7__2__0_left_grid_right_width_0_height_0_subtile_0__pin_ADDR_B1_i_0_),
		.right_width_0_height_1_subtile_0__pin_WDATA_A2_i_17_(cby_7__3__0_left_grid_right_width_0_height_1_subtile_0__pin_WDATA_A2_i_17_),
		.right_width_0_height_1_subtile_0__pin_ADDR_A2_i_1_(cby_7__3__0_left_grid_right_width_0_height_1_subtile_0__pin_ADDR_A2_i_1_),
		.right_width_0_height_1_subtile_0__pin_REN_A1_i_0_(cby_7__3__0_left_grid_right_width_0_height_1_subtile_0__pin_REN_A1_i_0_),
		.right_width_0_height_1_subtile_0__pin_REN_A2_i_0_(cby_7__3__0_left_grid_right_width_0_height_1_subtile_0__pin_REN_A2_i_0_),
		.right_width_0_height_1_subtile_0__pin_WEN_A2_i_0_(cby_7__3__0_left_grid_right_width_0_height_1_subtile_0__pin_WEN_A2_i_0_),
		.right_width_0_height_1_subtile_0__pin_BE_A2_i_0_(cby_7__3__0_left_grid_right_width_0_height_1_subtile_0__pin_BE_A2_i_0_),
		.right_width_0_height_1_subtile_0__pin_BE_A2_i_1_(cby_7__3__0_left_grid_right_width_0_height_1_subtile_0__pin_BE_A2_i_1_),
		.right_width_0_height_1_subtile_0__pin_WDATA_B1_i_0_(cby_7__3__0_left_grid_right_width_0_height_1_subtile_0__pin_WDATA_B1_i_0_),
		.right_width_0_height_1_subtile_0__pin_ADDR_B1_i_2_(cby_7__3__0_left_grid_right_width_0_height_1_subtile_0__pin_ADDR_B1_i_2_),
		.right_width_0_height_1_subtile_0__pin_ADDR_B1_i_3_(cby_7__3__0_left_grid_right_width_0_height_1_subtile_0__pin_ADDR_B1_i_3_),
		.right_width_0_height_1_subtile_0__pin_ADDR_B1_i_4_(cby_7__3__0_left_grid_right_width_0_height_1_subtile_0__pin_ADDR_B1_i_4_),
		.right_width_0_height_1_subtile_0__pin_ADDR_B1_i_5_(cby_7__3__0_left_grid_right_width_0_height_1_subtile_0__pin_ADDR_B1_i_5_),
		.right_width_0_height_1_subtile_0__pin_ADDR_B1_i_6_(cby_7__3__0_left_grid_right_width_0_height_1_subtile_0__pin_ADDR_B1_i_6_),
		.right_width_0_height_1_subtile_0__pin_ADDR_B1_i_7_(cby_7__3__0_left_grid_right_width_0_height_1_subtile_0__pin_ADDR_B1_i_7_),
		.right_width_0_height_1_subtile_0__pin_ADDR_B1_i_8_(cby_7__3__0_left_grid_right_width_0_height_1_subtile_0__pin_ADDR_B1_i_8_),
		.right_width_0_height_1_subtile_0__pin_ADDR_B1_i_9_(cby_7__3__0_left_grid_right_width_0_height_1_subtile_0__pin_ADDR_B1_i_9_),
		.right_width_0_height_1_subtile_0__pin_ADDR_B1_i_10_(cby_7__3__0_left_grid_right_width_0_height_1_subtile_0__pin_ADDR_B1_i_10_),
		.right_width_0_height_1_subtile_0__pin_ADDR_B1_i_11_(cby_7__3__0_left_grid_right_width_0_height_1_subtile_0__pin_ADDR_B1_i_11_),
		.right_width_0_height_1_subtile_0__pin_ADDR_B1_i_12_(cby_7__3__0_left_grid_right_width_0_height_1_subtile_0__pin_ADDR_B1_i_12_),
		.right_width_0_height_1_subtile_0__pin_ADDR_B1_i_13_(cby_7__3__0_left_grid_right_width_0_height_1_subtile_0__pin_ADDR_B1_i_13_),
		.right_width_0_height_1_subtile_0__pin_ADDR_B1_i_14_(cby_7__3__0_left_grid_right_width_0_height_1_subtile_0__pin_ADDR_B1_i_14_),
		.right_width_0_height_1_subtile_0__pin_FLUSH2_i_0_(cby_7__3__0_left_grid_right_width_0_height_1_subtile_0__pin_FLUSH2_i_0_),
		.right_width_0_height_2_subtile_0__pin_WDATA_A2_i_9_(cby_7__4__0_left_grid_right_width_0_height_2_subtile_0__pin_WDATA_A2_i_9_),
		.right_width_0_height_2_subtile_0__pin_WDATA_A2_i_10_(cby_7__4__0_left_grid_right_width_0_height_2_subtile_0__pin_WDATA_A2_i_10_),
		.right_width_0_height_2_subtile_0__pin_WDATA_A2_i_11_(cby_7__4__0_left_grid_right_width_0_height_2_subtile_0__pin_WDATA_A2_i_11_),
		.right_width_0_height_2_subtile_0__pin_WDATA_A2_i_12_(cby_7__4__0_left_grid_right_width_0_height_2_subtile_0__pin_WDATA_A2_i_12_),
		.right_width_0_height_2_subtile_0__pin_WDATA_A2_i_13_(cby_7__4__0_left_grid_right_width_0_height_2_subtile_0__pin_WDATA_A2_i_13_),
		.right_width_0_height_2_subtile_0__pin_WDATA_A2_i_14_(cby_7__4__0_left_grid_right_width_0_height_2_subtile_0__pin_WDATA_A2_i_14_),
		.right_width_0_height_2_subtile_0__pin_WDATA_A2_i_15_(cby_7__4__0_left_grid_right_width_0_height_2_subtile_0__pin_WDATA_A2_i_15_),
		.right_width_0_height_2_subtile_0__pin_WDATA_A2_i_16_(cby_7__4__0_left_grid_right_width_0_height_2_subtile_0__pin_WDATA_A2_i_16_),
		.right_width_0_height_2_subtile_0__pin_ADDR_A2_i_0_(cby_7__4__0_left_grid_right_width_0_height_2_subtile_0__pin_ADDR_A2_i_0_),
		.right_width_0_height_2_subtile_0__pin_ADDR_A2_i_2_(cby_7__4__0_left_grid_right_width_0_height_2_subtile_0__pin_ADDR_A2_i_2_),
		.right_width_0_height_2_subtile_0__pin_ADDR_A2_i_3_(cby_7__4__0_left_grid_right_width_0_height_2_subtile_0__pin_ADDR_A2_i_3_),
		.right_width_0_height_2_subtile_0__pin_ADDR_A2_i_4_(cby_7__4__0_left_grid_right_width_0_height_2_subtile_0__pin_ADDR_A2_i_4_),
		.right_width_0_height_2_subtile_0__pin_ADDR_A2_i_5_(cby_7__4__0_left_grid_right_width_0_height_2_subtile_0__pin_ADDR_A2_i_5_),
		.right_width_0_height_2_subtile_0__pin_ADDR_A2_i_6_(cby_7__4__0_left_grid_right_width_0_height_2_subtile_0__pin_ADDR_A2_i_6_),
		.right_width_0_height_2_subtile_0__pin_ADDR_A2_i_7_(cby_7__4__0_left_grid_right_width_0_height_2_subtile_0__pin_ADDR_A2_i_7_),
		.right_width_0_height_2_subtile_0__pin_ADDR_A2_i_8_(cby_7__4__0_left_grid_right_width_0_height_2_subtile_0__pin_ADDR_A2_i_8_),
		.right_width_0_height_2_subtile_0__pin_ADDR_A2_i_9_(cby_7__4__0_left_grid_right_width_0_height_2_subtile_0__pin_ADDR_A2_i_9_),
		.right_width_0_height_2_subtile_0__pin_ADDR_A2_i_10_(cby_7__4__0_left_grid_right_width_0_height_2_subtile_0__pin_ADDR_A2_i_10_),
		.right_width_0_height_2_subtile_0__pin_ADDR_A2_i_11_(cby_7__4__0_left_grid_right_width_0_height_2_subtile_0__pin_ADDR_A2_i_11_),
		.right_width_0_height_2_subtile_0__pin_ADDR_A2_i_12_(cby_7__4__0_left_grid_right_width_0_height_2_subtile_0__pin_ADDR_A2_i_12_),
		.right_width_0_height_2_subtile_0__pin_ADDR_A2_i_13_(cby_7__4__0_left_grid_right_width_0_height_2_subtile_0__pin_ADDR_A2_i_13_),
		.right_width_0_height_2_subtile_0__pin_WEN_A1_i_0_(cby_7__4__0_left_grid_right_width_0_height_2_subtile_0__pin_WEN_A1_i_0_),
		.right_width_0_height_3_subtile_0__pin_WDATA_A1_i_7_(cby_7__5__0_left_grid_right_width_0_height_3_subtile_0__pin_WDATA_A1_i_7_),
		.right_width_0_height_3_subtile_0__pin_WDATA_A1_i_8_(cby_7__5__0_left_grid_right_width_0_height_3_subtile_0__pin_WDATA_A1_i_8_),
		.right_width_0_height_3_subtile_0__pin_WDATA_A1_i_9_(cby_7__5__0_left_grid_right_width_0_height_3_subtile_0__pin_WDATA_A1_i_9_),
		.right_width_0_height_3_subtile_0__pin_WDATA_A1_i_10_(cby_7__5__0_left_grid_right_width_0_height_3_subtile_0__pin_WDATA_A1_i_10_),
		.right_width_0_height_3_subtile_0__pin_WDATA_A1_i_11_(cby_7__5__0_left_grid_right_width_0_height_3_subtile_0__pin_WDATA_A1_i_11_),
		.right_width_0_height_3_subtile_0__pin_WDATA_A1_i_12_(cby_7__5__0_left_grid_right_width_0_height_3_subtile_0__pin_WDATA_A1_i_12_),
		.right_width_0_height_3_subtile_0__pin_WDATA_A1_i_13_(cby_7__5__0_left_grid_right_width_0_height_3_subtile_0__pin_WDATA_A1_i_13_),
		.right_width_0_height_3_subtile_0__pin_WDATA_A1_i_14_(cby_7__5__0_left_grid_right_width_0_height_3_subtile_0__pin_WDATA_A1_i_14_),
		.right_width_0_height_3_subtile_0__pin_WDATA_A1_i_15_(cby_7__5__0_left_grid_right_width_0_height_3_subtile_0__pin_WDATA_A1_i_15_),
		.right_width_0_height_3_subtile_0__pin_WDATA_A1_i_16_(cby_7__5__0_left_grid_right_width_0_height_3_subtile_0__pin_WDATA_A1_i_16_),
		.right_width_0_height_3_subtile_0__pin_WDATA_A1_i_17_(cby_7__5__0_left_grid_right_width_0_height_3_subtile_0__pin_WDATA_A1_i_17_),
		.right_width_0_height_3_subtile_0__pin_ADDR_A1_i_0_(cby_7__5__0_left_grid_right_width_0_height_3_subtile_0__pin_ADDR_A1_i_0_),
		.right_width_0_height_3_subtile_0__pin_ADDR_A1_i_1_(cby_7__5__0_left_grid_right_width_0_height_3_subtile_0__pin_ADDR_A1_i_1_),
		.right_width_0_height_3_subtile_0__pin_BE_A1_i_0_(cby_7__5__0_left_grid_right_width_0_height_3_subtile_0__pin_BE_A1_i_0_),
		.right_width_0_height_3_subtile_0__pin_BE_A1_i_1_(cby_7__5__0_left_grid_right_width_0_height_3_subtile_0__pin_BE_A1_i_1_),
		.right_width_0_height_3_subtile_0__pin_REN_B2_i_0_(cby_7__5__0_left_grid_right_width_0_height_3_subtile_0__pin_REN_B2_i_0_),
		.right_width_0_height_3_subtile_0__pin_WEN_B2_i_0_(cby_7__5__0_left_grid_right_width_0_height_3_subtile_0__pin_WEN_B2_i_0_),
		.right_width_0_height_3_subtile_0__pin_BE_B1_i_0_(cby_7__5__0_left_grid_right_width_0_height_3_subtile_0__pin_BE_B1_i_0_),
		.right_width_0_height_3_subtile_0__pin_BE_B1_i_1_(cby_7__5__0_left_grid_right_width_0_height_3_subtile_0__pin_BE_B1_i_1_),
		.right_width_0_height_3_subtile_0__pin_BE_B2_i_0_(cby_7__5__0_left_grid_right_width_0_height_3_subtile_0__pin_BE_B2_i_0_),
		.right_width_0_height_3_subtile_0__pin_BE_B2_i_1_(cby_7__5__0_left_grid_right_width_0_height_3_subtile_0__pin_BE_B2_i_1_),
		.right_width_0_height_3_subtile_0__pin_FLUSH1_i_0_(cby_7__5__0_left_grid_right_width_0_height_3_subtile_0__pin_FLUSH1_i_0_),
		.right_width_0_height_4_subtile_0__pin_WDATA_A2_i_0_(cby_7__6__0_left_grid_right_width_0_height_4_subtile_0__pin_WDATA_A2_i_0_),
		.right_width_0_height_4_subtile_0__pin_WDATA_A2_i_1_(cby_7__6__0_left_grid_right_width_0_height_4_subtile_0__pin_WDATA_A2_i_1_),
		.right_width_0_height_4_subtile_0__pin_WDATA_A2_i_2_(cby_7__6__0_left_grid_right_width_0_height_4_subtile_0__pin_WDATA_A2_i_2_),
		.right_width_0_height_4_subtile_0__pin_WDATA_A2_i_3_(cby_7__6__0_left_grid_right_width_0_height_4_subtile_0__pin_WDATA_A2_i_3_),
		.right_width_0_height_4_subtile_0__pin_WDATA_A2_i_4_(cby_7__6__0_left_grid_right_width_0_height_4_subtile_0__pin_WDATA_A2_i_4_),
		.right_width_0_height_4_subtile_0__pin_WDATA_A2_i_5_(cby_7__6__0_left_grid_right_width_0_height_4_subtile_0__pin_WDATA_A2_i_5_),
		.right_width_0_height_4_subtile_0__pin_WDATA_A2_i_6_(cby_7__6__0_left_grid_right_width_0_height_4_subtile_0__pin_WDATA_A2_i_6_),
		.right_width_0_height_4_subtile_0__pin_WDATA_A2_i_7_(cby_7__6__0_left_grid_right_width_0_height_4_subtile_0__pin_WDATA_A2_i_7_),
		.right_width_0_height_4_subtile_0__pin_WDATA_A2_i_8_(cby_7__6__0_left_grid_right_width_0_height_4_subtile_0__pin_WDATA_A2_i_8_),
		.right_width_0_height_4_subtile_0__pin_WDATA_B2_i_17_(cby_7__6__0_left_grid_right_width_0_height_4_subtile_0__pin_WDATA_B2_i_17_),
		.right_width_0_height_4_subtile_0__pin_ADDR_B2_i_1_(cby_7__6__0_left_grid_right_width_0_height_4_subtile_0__pin_ADDR_B2_i_1_),
		.right_width_0_height_4_subtile_0__pin_ADDR_B2_i_4_(cby_7__6__0_left_grid_right_width_0_height_4_subtile_0__pin_ADDR_B2_i_4_),
		.right_width_0_height_4_subtile_0__pin_ADDR_B2_i_5_(cby_7__6__0_left_grid_right_width_0_height_4_subtile_0__pin_ADDR_B2_i_5_),
		.right_width_0_height_4_subtile_0__pin_ADDR_B2_i_6_(cby_7__6__0_left_grid_right_width_0_height_4_subtile_0__pin_ADDR_B2_i_6_),
		.right_width_0_height_4_subtile_0__pin_ADDR_B2_i_7_(cby_7__6__0_left_grid_right_width_0_height_4_subtile_0__pin_ADDR_B2_i_7_),
		.right_width_0_height_4_subtile_0__pin_ADDR_B2_i_8_(cby_7__6__0_left_grid_right_width_0_height_4_subtile_0__pin_ADDR_B2_i_8_),
		.right_width_0_height_4_subtile_0__pin_ADDR_B2_i_9_(cby_7__6__0_left_grid_right_width_0_height_4_subtile_0__pin_ADDR_B2_i_9_),
		.right_width_0_height_4_subtile_0__pin_ADDR_B2_i_10_(cby_7__6__0_left_grid_right_width_0_height_4_subtile_0__pin_ADDR_B2_i_10_),
		.right_width_0_height_4_subtile_0__pin_ADDR_B2_i_11_(cby_7__6__0_left_grid_right_width_0_height_4_subtile_0__pin_ADDR_B2_i_11_),
		.right_width_0_height_4_subtile_0__pin_ADDR_B2_i_12_(cby_7__6__0_left_grid_right_width_0_height_4_subtile_0__pin_ADDR_B2_i_12_),
		.right_width_0_height_4_subtile_0__pin_ADDR_B2_i_13_(cby_7__6__0_left_grid_right_width_0_height_4_subtile_0__pin_ADDR_B2_i_13_),
		.right_width_0_height_4_subtile_0__pin_WEN_B1_i_0_(cby_7__6__0_left_grid_right_width_0_height_4_subtile_0__pin_WEN_B1_i_0_),
		.right_width_0_height_5_subtile_0__pin_WDATA_B2_i_0_(cby_7__7__0_left_grid_right_width_0_height_5_subtile_0__pin_WDATA_B2_i_0_),
		.right_width_0_height_5_subtile_0__pin_WDATA_B2_i_1_(cby_7__7__0_left_grid_right_width_0_height_5_subtile_0__pin_WDATA_B2_i_1_),
		.right_width_0_height_5_subtile_0__pin_WDATA_B2_i_2_(cby_7__7__0_left_grid_right_width_0_height_5_subtile_0__pin_WDATA_B2_i_2_),
		.right_width_0_height_5_subtile_0__pin_WDATA_B2_i_3_(cby_7__7__0_left_grid_right_width_0_height_5_subtile_0__pin_WDATA_B2_i_3_),
		.right_width_0_height_5_subtile_0__pin_WDATA_B2_i_4_(cby_7__7__0_left_grid_right_width_0_height_5_subtile_0__pin_WDATA_B2_i_4_),
		.right_width_0_height_5_subtile_0__pin_WDATA_B2_i_5_(cby_7__7__0_left_grid_right_width_0_height_5_subtile_0__pin_WDATA_B2_i_5_),
		.right_width_0_height_5_subtile_0__pin_WDATA_B2_i_6_(cby_7__7__0_left_grid_right_width_0_height_5_subtile_0__pin_WDATA_B2_i_6_),
		.right_width_0_height_5_subtile_0__pin_WDATA_B2_i_7_(cby_7__7__0_left_grid_right_width_0_height_5_subtile_0__pin_WDATA_B2_i_7_),
		.right_width_0_height_5_subtile_0__pin_WDATA_B2_i_8_(cby_7__7__0_left_grid_right_width_0_height_5_subtile_0__pin_WDATA_B2_i_8_),
		.right_width_0_height_5_subtile_0__pin_WDATA_B2_i_9_(cby_7__7__0_left_grid_right_width_0_height_5_subtile_0__pin_WDATA_B2_i_9_),
		.right_width_0_height_5_subtile_0__pin_WDATA_B2_i_10_(cby_7__7__0_left_grid_right_width_0_height_5_subtile_0__pin_WDATA_B2_i_10_),
		.right_width_0_height_5_subtile_0__pin_WDATA_B2_i_11_(cby_7__7__0_left_grid_right_width_0_height_5_subtile_0__pin_WDATA_B2_i_11_),
		.right_width_0_height_5_subtile_0__pin_WDATA_B2_i_12_(cby_7__7__0_left_grid_right_width_0_height_5_subtile_0__pin_WDATA_B2_i_12_),
		.right_width_0_height_5_subtile_0__pin_WDATA_B2_i_13_(cby_7__7__0_left_grid_right_width_0_height_5_subtile_0__pin_WDATA_B2_i_13_),
		.right_width_0_height_5_subtile_0__pin_WDATA_B2_i_14_(cby_7__7__0_left_grid_right_width_0_height_5_subtile_0__pin_WDATA_B2_i_14_),
		.right_width_0_height_5_subtile_0__pin_WDATA_B2_i_15_(cby_7__7__0_left_grid_right_width_0_height_5_subtile_0__pin_WDATA_B2_i_15_),
		.right_width_0_height_5_subtile_0__pin_WDATA_B2_i_16_(cby_7__7__0_left_grid_right_width_0_height_5_subtile_0__pin_WDATA_B2_i_16_),
		.right_width_0_height_5_subtile_0__pin_ADDR_B2_i_0_(cby_7__7__0_left_grid_right_width_0_height_5_subtile_0__pin_ADDR_B2_i_0_),
		.right_width_0_height_5_subtile_0__pin_ADDR_B2_i_2_(cby_7__7__0_left_grid_right_width_0_height_5_subtile_0__pin_ADDR_B2_i_2_),
		.right_width_0_height_5_subtile_0__pin_ADDR_B2_i_3_(cby_7__7__0_left_grid_right_width_0_height_5_subtile_0__pin_ADDR_B2_i_3_),
		.right_width_0_height_5_subtile_0__pin_REN_B1_i_0_(cby_7__7__0_left_grid_right_width_0_height_5_subtile_0__pin_REN_B1_i_0_),
		.bottom_width_0_height_0_subtile_0__pin_WDATA_A1_i_0_(cbx_7__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_WDATA_A1_i_0_),
		.bottom_width_0_height_0_subtile_0__pin_WDATA_A1_i_1_(cbx_7__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_WDATA_A1_i_1_),
		.bottom_width_0_height_0_subtile_0__pin_WDATA_A1_i_2_(cbx_7__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_WDATA_A1_i_2_),
		.bottom_width_0_height_0_subtile_0__pin_WDATA_A1_i_3_(cbx_7__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_WDATA_A1_i_3_),
		.bottom_width_0_height_0_subtile_0__pin_WDATA_A1_i_4_(cbx_7__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_WDATA_A1_i_4_),
		.bottom_width_0_height_0_subtile_0__pin_WDATA_A1_i_5_(cbx_7__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_WDATA_A1_i_5_),
		.bottom_width_0_height_0_subtile_0__pin_WDATA_A1_i_6_(cbx_7__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_WDATA_A1_i_6_),
		.bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_6_(cbx_7__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_6_),
		.bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_7_(cbx_7__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_7_),
		.bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_8_(cbx_7__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_8_),
		.bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_9_(cbx_7__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_9_),
		.bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_10_(cbx_7__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_10_),
		.bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_11_(cbx_7__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_11_),
		.bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_12_(cbx_7__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_12_),
		.bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_13_(cbx_7__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_13_),
		.bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_14_(cbx_7__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_14_),
		.bottom_width_0_height_0_subtile_0__pin_WDATA_B1_i_17_(cbx_7__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_WDATA_B1_i_17_),
		.bottom_width_0_height_0_subtile_0__pin_ADDR_B1_i_1_(cbx_7__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ADDR_B1_i_1_),
		.left_width_0_height_0_subtile_0__pin_RAM_ID_i_0_(grid_bram_7__2__undriven_left_width_0_height_0_subtile_0__pin_RAM_ID_i_0_),
		.left_width_0_height_0_subtile_0__pin_RAM_ID_i_1_(grid_bram_7__2__undriven_left_width_0_height_0_subtile_0__pin_RAM_ID_i_1_),
		.left_width_0_height_0_subtile_0__pin_RAM_ID_i_2_(grid_bram_7__2__undriven_left_width_0_height_0_subtile_0__pin_RAM_ID_i_2_),
		.left_width_0_height_0_subtile_0__pin_RAM_ID_i_3_(grid_bram_7__2__undriven_left_width_0_height_0_subtile_0__pin_RAM_ID_i_3_),
		.left_width_0_height_0_subtile_0__pin_RAM_ID_i_4_(grid_bram_7__2__undriven_left_width_0_height_0_subtile_0__pin_RAM_ID_i_4_),
		.left_width_0_height_0_subtile_0__pin_RAM_ID_i_5_(grid_bram_7__2__undriven_left_width_0_height_0_subtile_0__pin_RAM_ID_i_5_),
		.left_width_0_height_0_subtile_0__pin_RAM_ID_i_6_(grid_bram_7__2__undriven_left_width_0_height_0_subtile_0__pin_RAM_ID_i_6_),
		.left_width_0_height_0_subtile_0__pin_RAM_ID_i_7_(grid_bram_7__2__undriven_left_width_0_height_0_subtile_0__pin_RAM_ID_i_7_),
		.left_width_0_height_0_subtile_0__pin_RAM_ID_i_8_(grid_bram_7__2__undriven_left_width_0_height_0_subtile_0__pin_RAM_ID_i_8_),
		.left_width_0_height_0_subtile_0__pin_RAM_ID_i_9_(grid_bram_7__2__undriven_left_width_0_height_0_subtile_0__pin_RAM_ID_i_9_),
		.left_width_0_height_0_subtile_0__pin_RAM_ID_i_10_(grid_bram_7__2__undriven_left_width_0_height_0_subtile_0__pin_RAM_ID_i_10_),
		.left_width_0_height_0_subtile_0__pin_RAM_ID_i_11_(grid_bram_7__2__undriven_left_width_0_height_0_subtile_0__pin_RAM_ID_i_11_),
		.left_width_0_height_0_subtile_0__pin_RAM_ID_i_12_(grid_bram_7__2__undriven_left_width_0_height_0_subtile_0__pin_RAM_ID_i_12_),
		.left_width_0_height_0_subtile_0__pin_RAM_ID_i_13_(grid_bram_7__2__undriven_left_width_0_height_0_subtile_0__pin_RAM_ID_i_13_),
		.left_width_0_height_0_subtile_0__pin_RAM_ID_i_14_(grid_bram_7__2__undriven_left_width_0_height_0_subtile_0__pin_RAM_ID_i_14_),
		.left_width_0_height_0_subtile_0__pin_RAM_ID_i_15_(grid_bram_7__2__undriven_left_width_0_height_0_subtile_0__pin_RAM_ID_i_15_),
		.left_width_0_height_0_subtile_0__pin_RAM_ID_i_16_(grid_bram_7__2__undriven_left_width_0_height_0_subtile_0__pin_RAM_ID_i_16_),
		.left_width_0_height_0_subtile_0__pin_RAM_ID_i_17_(grid_bram_7__2__undriven_left_width_0_height_0_subtile_0__pin_RAM_ID_i_17_),
		.left_width_0_height_0_subtile_0__pin_RAM_ID_i_18_(grid_bram_7__2__undriven_left_width_0_height_0_subtile_0__pin_RAM_ID_i_18_),
		.left_width_0_height_0_subtile_0__pin_RAM_ID_i_19_(grid_bram_7__2__undriven_left_width_0_height_0_subtile_0__pin_RAM_ID_i_19_),
		.left_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.ccff_head(cby_7__2__0_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_RDATA_A1_o_0_(grid_bram_0_right_width_0_height_0_subtile_0__pin_RDATA_A1_o_0_),
		.right_width_0_height_0_subtile_0__pin_RDATA_A1_o_1_(grid_bram_0_right_width_0_height_0_subtile_0__pin_RDATA_A1_o_1_),
		.right_width_0_height_0_subtile_0__pin_RDATA_A1_o_2_(grid_bram_0_right_width_0_height_0_subtile_0__pin_RDATA_A1_o_2_),
		.right_width_0_height_0_subtile_0__pin_RDATA_A1_o_3_(grid_bram_0_right_width_0_height_0_subtile_0__pin_RDATA_A1_o_3_),
		.right_width_0_height_0_subtile_0__pin_RDATA_A1_o_4_(grid_bram_0_right_width_0_height_0_subtile_0__pin_RDATA_A1_o_4_),
		.right_width_0_height_0_subtile_0__pin_RDATA_A1_o_5_(grid_bram_0_right_width_0_height_0_subtile_0__pin_RDATA_A1_o_5_),
		.right_width_0_height_0_subtile_0__pin_RDATA_B1_o_0_(grid_bram_0_right_width_0_height_0_subtile_0__pin_RDATA_B1_o_0_),
		.right_width_0_height_0_subtile_0__pin_RDATA_B1_o_1_(grid_bram_0_right_width_0_height_0_subtile_0__pin_RDATA_B1_o_1_),
		.right_width_0_height_0_subtile_0__pin_RDATA_B1_o_2_(grid_bram_0_right_width_0_height_0_subtile_0__pin_RDATA_B1_o_2_),
		.right_width_0_height_0_subtile_0__pin_RDATA_B1_o_3_(grid_bram_0_right_width_0_height_0_subtile_0__pin_RDATA_B1_o_3_),
		.right_width_0_height_0_subtile_0__pin_RDATA_B1_o_4_(grid_bram_0_right_width_0_height_0_subtile_0__pin_RDATA_B1_o_4_),
		.right_width_0_height_0_subtile_0__pin_RDATA_B1_o_5_(grid_bram_0_right_width_0_height_0_subtile_0__pin_RDATA_B1_o_5_),
		.right_width_0_height_1_subtile_0__pin_RDATA_A1_o_6_(grid_bram_0_right_width_0_height_1_subtile_0__pin_RDATA_A1_o_6_),
		.right_width_0_height_1_subtile_0__pin_RDATA_A1_o_7_(grid_bram_0_right_width_0_height_1_subtile_0__pin_RDATA_A1_o_7_),
		.right_width_0_height_1_subtile_0__pin_RDATA_A1_o_8_(grid_bram_0_right_width_0_height_1_subtile_0__pin_RDATA_A1_o_8_),
		.right_width_0_height_1_subtile_0__pin_RDATA_A1_o_9_(grid_bram_0_right_width_0_height_1_subtile_0__pin_RDATA_A1_o_9_),
		.right_width_0_height_1_subtile_0__pin_RDATA_A1_o_10_(grid_bram_0_right_width_0_height_1_subtile_0__pin_RDATA_A1_o_10_),
		.right_width_0_height_1_subtile_0__pin_RDATA_A1_o_11_(grid_bram_0_right_width_0_height_1_subtile_0__pin_RDATA_A1_o_11_),
		.right_width_0_height_1_subtile_0__pin_RDATA_B1_o_6_(grid_bram_0_right_width_0_height_1_subtile_0__pin_RDATA_B1_o_6_),
		.right_width_0_height_1_subtile_0__pin_RDATA_B1_o_7_(grid_bram_0_right_width_0_height_1_subtile_0__pin_RDATA_B1_o_7_),
		.right_width_0_height_1_subtile_0__pin_RDATA_B1_o_8_(grid_bram_0_right_width_0_height_1_subtile_0__pin_RDATA_B1_o_8_),
		.right_width_0_height_1_subtile_0__pin_RDATA_B1_o_9_(grid_bram_0_right_width_0_height_1_subtile_0__pin_RDATA_B1_o_9_),
		.right_width_0_height_1_subtile_0__pin_RDATA_B1_o_10_(grid_bram_0_right_width_0_height_1_subtile_0__pin_RDATA_B1_o_10_),
		.right_width_0_height_1_subtile_0__pin_RDATA_B1_o_11_(grid_bram_0_right_width_0_height_1_subtile_0__pin_RDATA_B1_o_11_),
		.right_width_0_height_2_subtile_0__pin_RDATA_A1_o_12_(grid_bram_0_right_width_0_height_2_subtile_0__pin_RDATA_A1_o_12_),
		.right_width_0_height_2_subtile_0__pin_RDATA_A1_o_13_(grid_bram_0_right_width_0_height_2_subtile_0__pin_RDATA_A1_o_13_),
		.right_width_0_height_2_subtile_0__pin_RDATA_A1_o_14_(grid_bram_0_right_width_0_height_2_subtile_0__pin_RDATA_A1_o_14_),
		.right_width_0_height_2_subtile_0__pin_RDATA_A1_o_15_(grid_bram_0_right_width_0_height_2_subtile_0__pin_RDATA_A1_o_15_),
		.right_width_0_height_2_subtile_0__pin_RDATA_A1_o_16_(grid_bram_0_right_width_0_height_2_subtile_0__pin_RDATA_A1_o_16_),
		.right_width_0_height_2_subtile_0__pin_RDATA_A1_o_17_(grid_bram_0_right_width_0_height_2_subtile_0__pin_RDATA_A1_o_17_),
		.right_width_0_height_2_subtile_0__pin_RDATA_B1_o_12_(grid_bram_0_right_width_0_height_2_subtile_0__pin_RDATA_B1_o_12_),
		.right_width_0_height_2_subtile_0__pin_RDATA_B1_o_13_(grid_bram_0_right_width_0_height_2_subtile_0__pin_RDATA_B1_o_13_),
		.right_width_0_height_2_subtile_0__pin_RDATA_B1_o_14_(grid_bram_0_right_width_0_height_2_subtile_0__pin_RDATA_B1_o_14_),
		.right_width_0_height_2_subtile_0__pin_RDATA_B1_o_15_(grid_bram_0_right_width_0_height_2_subtile_0__pin_RDATA_B1_o_15_),
		.right_width_0_height_2_subtile_0__pin_RDATA_B1_o_16_(grid_bram_0_right_width_0_height_2_subtile_0__pin_RDATA_B1_o_16_),
		.right_width_0_height_2_subtile_0__pin_RDATA_B1_o_17_(grid_bram_0_right_width_0_height_2_subtile_0__pin_RDATA_B1_o_17_),
		.right_width_0_height_3_subtile_0__pin_RDATA_A2_o_0_(grid_bram_0_right_width_0_height_3_subtile_0__pin_RDATA_A2_o_0_),
		.right_width_0_height_3_subtile_0__pin_RDATA_A2_o_1_(grid_bram_0_right_width_0_height_3_subtile_0__pin_RDATA_A2_o_1_),
		.right_width_0_height_3_subtile_0__pin_RDATA_A2_o_2_(grid_bram_0_right_width_0_height_3_subtile_0__pin_RDATA_A2_o_2_),
		.right_width_0_height_3_subtile_0__pin_RDATA_A2_o_3_(grid_bram_0_right_width_0_height_3_subtile_0__pin_RDATA_A2_o_3_),
		.right_width_0_height_3_subtile_0__pin_RDATA_A2_o_4_(grid_bram_0_right_width_0_height_3_subtile_0__pin_RDATA_A2_o_4_),
		.right_width_0_height_3_subtile_0__pin_RDATA_A2_o_5_(grid_bram_0_right_width_0_height_3_subtile_0__pin_RDATA_A2_o_5_),
		.right_width_0_height_3_subtile_0__pin_RDATA_B2_o_0_(grid_bram_0_right_width_0_height_3_subtile_0__pin_RDATA_B2_o_0_),
		.right_width_0_height_3_subtile_0__pin_RDATA_B2_o_1_(grid_bram_0_right_width_0_height_3_subtile_0__pin_RDATA_B2_o_1_),
		.right_width_0_height_3_subtile_0__pin_RDATA_B2_o_2_(grid_bram_0_right_width_0_height_3_subtile_0__pin_RDATA_B2_o_2_),
		.right_width_0_height_3_subtile_0__pin_RDATA_B2_o_3_(grid_bram_0_right_width_0_height_3_subtile_0__pin_RDATA_B2_o_3_),
		.right_width_0_height_3_subtile_0__pin_RDATA_B2_o_4_(grid_bram_0_right_width_0_height_3_subtile_0__pin_RDATA_B2_o_4_),
		.right_width_0_height_3_subtile_0__pin_RDATA_B2_o_5_(grid_bram_0_right_width_0_height_3_subtile_0__pin_RDATA_B2_o_5_),
		.right_width_0_height_4_subtile_0__pin_RDATA_A2_o_6_(grid_bram_0_right_width_0_height_4_subtile_0__pin_RDATA_A2_o_6_),
		.right_width_0_height_4_subtile_0__pin_RDATA_A2_o_7_(grid_bram_0_right_width_0_height_4_subtile_0__pin_RDATA_A2_o_7_),
		.right_width_0_height_4_subtile_0__pin_RDATA_A2_o_8_(grid_bram_0_right_width_0_height_4_subtile_0__pin_RDATA_A2_o_8_),
		.right_width_0_height_4_subtile_0__pin_RDATA_A2_o_9_(grid_bram_0_right_width_0_height_4_subtile_0__pin_RDATA_A2_o_9_),
		.right_width_0_height_4_subtile_0__pin_RDATA_A2_o_10_(grid_bram_0_right_width_0_height_4_subtile_0__pin_RDATA_A2_o_10_),
		.right_width_0_height_4_subtile_0__pin_RDATA_A2_o_11_(grid_bram_0_right_width_0_height_4_subtile_0__pin_RDATA_A2_o_11_),
		.right_width_0_height_4_subtile_0__pin_RDATA_B2_o_6_(grid_bram_0_right_width_0_height_4_subtile_0__pin_RDATA_B2_o_6_),
		.right_width_0_height_4_subtile_0__pin_RDATA_B2_o_7_(grid_bram_0_right_width_0_height_4_subtile_0__pin_RDATA_B2_o_7_),
		.right_width_0_height_4_subtile_0__pin_RDATA_B2_o_8_(grid_bram_0_right_width_0_height_4_subtile_0__pin_RDATA_B2_o_8_),
		.right_width_0_height_4_subtile_0__pin_RDATA_B2_o_9_(grid_bram_0_right_width_0_height_4_subtile_0__pin_RDATA_B2_o_9_),
		.right_width_0_height_4_subtile_0__pin_RDATA_B2_o_10_(grid_bram_0_right_width_0_height_4_subtile_0__pin_RDATA_B2_o_10_),
		.right_width_0_height_4_subtile_0__pin_RDATA_B2_o_11_(grid_bram_0_right_width_0_height_4_subtile_0__pin_RDATA_B2_o_11_),
		.right_width_0_height_5_subtile_0__pin_RDATA_A2_o_12_(grid_bram_0_right_width_0_height_5_subtile_0__pin_RDATA_A2_o_12_),
		.right_width_0_height_5_subtile_0__pin_RDATA_A2_o_13_(grid_bram_0_right_width_0_height_5_subtile_0__pin_RDATA_A2_o_13_),
		.right_width_0_height_5_subtile_0__pin_RDATA_A2_o_14_(grid_bram_0_right_width_0_height_5_subtile_0__pin_RDATA_A2_o_14_),
		.right_width_0_height_5_subtile_0__pin_RDATA_A2_o_15_(grid_bram_0_right_width_0_height_5_subtile_0__pin_RDATA_A2_o_15_),
		.right_width_0_height_5_subtile_0__pin_RDATA_A2_o_16_(grid_bram_0_right_width_0_height_5_subtile_0__pin_RDATA_A2_o_16_),
		.right_width_0_height_5_subtile_0__pin_RDATA_A2_o_17_(grid_bram_0_right_width_0_height_5_subtile_0__pin_RDATA_A2_o_17_),
		.right_width_0_height_5_subtile_0__pin_RDATA_B2_o_12_(grid_bram_0_right_width_0_height_5_subtile_0__pin_RDATA_B2_o_12_),
		.right_width_0_height_5_subtile_0__pin_RDATA_B2_o_13_(grid_bram_0_right_width_0_height_5_subtile_0__pin_RDATA_B2_o_13_),
		.right_width_0_height_5_subtile_0__pin_RDATA_B2_o_14_(grid_bram_0_right_width_0_height_5_subtile_0__pin_RDATA_B2_o_14_),
		.right_width_0_height_5_subtile_0__pin_RDATA_B2_o_15_(grid_bram_0_right_width_0_height_5_subtile_0__pin_RDATA_B2_o_15_),
		.right_width_0_height_5_subtile_0__pin_RDATA_B2_o_16_(grid_bram_0_right_width_0_height_5_subtile_0__pin_RDATA_B2_o_16_),
		.right_width_0_height_5_subtile_0__pin_RDATA_B2_o_17_(grid_bram_0_right_width_0_height_5_subtile_0__pin_RDATA_B2_o_17_),
		.bottom_width_0_height_0_subtile_0__pin_PL_INIT_o_0_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_INIT_o_0_),
		.bottom_width_0_height_0_subtile_0__pin_PL_ENA_o_0_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_ENA_o_0_),
		.bottom_width_0_height_0_subtile_0__pin_PL_REN_o_0_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_REN_o_0_),
		.bottom_width_0_height_0_subtile_0__pin_PL_CLK_o_0_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_CLK_o_0_),
		.bottom_width_0_height_0_subtile_0__pin_PL_WEN_o_0_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_WEN_o_0_),
		.bottom_width_0_height_0_subtile_0__pin_PL_WEN_o_1_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_WEN_o_1_),
		.bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_0_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_0_),
		.bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_1_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_1_),
		.bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_2_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_2_),
		.bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_3_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_3_),
		.bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_4_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_4_),
		.bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_5_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_5_),
		.bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_6_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_6_),
		.bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_7_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_7_),
		.bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_8_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_8_),
		.bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_9_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_9_),
		.bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_10_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_10_),
		.bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_11_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_11_),
		.bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_12_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_12_),
		.bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_13_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_13_),
		.bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_14_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_14_),
		.bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_15_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_15_),
		.bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_16_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_16_),
		.bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_17_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_17_),
		.bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_18_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_18_),
		.bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_19_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_19_),
		.bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_20_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_20_),
		.bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_21_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_21_),
		.bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_22_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_22_),
		.bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_23_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_23_),
		.bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_24_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_24_),
		.bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_25_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_25_),
		.bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_26_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_26_),
		.bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_27_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_27_),
		.bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_28_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_28_),
		.bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_29_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_29_),
		.bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_30_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_30_),
		.bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_31_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_31_),
		.bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_0_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_0_),
		.bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_1_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_1_),
		.bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_2_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_2_),
		.bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_3_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_3_),
		.bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_4_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_4_),
		.bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_5_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_5_),
		.bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_6_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_6_),
		.bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_7_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_7_),
		.bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_8_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_8_),
		.bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_9_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_9_),
		.bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_10_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_10_),
		.bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_11_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_11_),
		.bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_12_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_12_),
		.bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_13_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_13_),
		.bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_14_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_14_),
		.bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_15_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_15_),
		.bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_16_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_16_),
		.bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_17_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_17_),
		.bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_18_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_18_),
		.bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_19_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_19_),
		.bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_20_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_20_),
		.bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_21_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_21_),
		.bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_22_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_22_),
		.bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_23_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_23_),
		.bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_24_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_24_),
		.bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_25_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_25_),
		.bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_26_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_26_),
		.bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_27_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_27_),
		.bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_28_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_28_),
		.bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_29_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_29_),
		.bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_30_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_30_),
		.bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_31_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_31_),
		.bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_32_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_32_),
		.bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_33_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_33_),
		.bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_34_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_34_),
		.bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_35_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_35_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_1_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_1_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_2_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_2_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_3_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_3_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_4_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_4_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_5_(grid_bram_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_5_),
		.ccff_tail(grid_bram_0_ccff_tail));

	grid_io_right grid_io_right_10__1_ (
		.test_en(test_en),
		.scan_mode(scan_mode),
		.scan_clk(scan_clk),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.CFG_DONE(CFG_DONE),
		.gfpga_pad_QL_PREIO_A2F(gfpga_pad_QL_PREIO_A2F[460:479]),
		.gfpga_pad_QL_PREIO_F2A(gfpga_pad_QL_PREIO_F2A[460:479]),
		.gfpga_pad_QL_PREIO_F2A_DEF0(gfpga_pad_QL_PREIO_F2A_DEF0[460:479]),
		.gfpga_pad_QL_PREIO_F2A_DEF1(gfpga_pad_QL_PREIO_F2A_DEF1[460:479]),
		.gfpga_pad_QL_PREIO_F2A_CLK(gfpga_pad_QL_PREIO_F2A_CLK[460:479]),
		.left_width_0_height_0_subtile_0__pin_f2a_i_0_(cby_9__1__0_right_grid_left_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_0__pin_sc_in_0_(grid_io_right_10__1__undriven_left_width_0_height_0_subtile_0__pin_sc_in_0_),
		.left_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_1__pin_f2a_i_0_(cby_9__1__0_right_grid_left_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_1__pin_sc_in_0_(grid_io_right_10__1__undriven_left_width_0_height_0_subtile_1__pin_sc_in_0_),
		.left_width_0_height_0_subtile_1__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_1__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_1__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_1__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_1__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_1__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_2__pin_f2a_i_0_(cby_9__1__0_right_grid_left_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_2__pin_sc_in_0_(grid_io_right_10__1__undriven_left_width_0_height_0_subtile_2__pin_sc_in_0_),
		.left_width_0_height_0_subtile_2__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_2__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_2__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_2__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_2__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_2__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_3__pin_f2a_i_0_(cby_9__1__0_right_grid_left_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_3__pin_sc_in_0_(grid_io_right_10__1__undriven_left_width_0_height_0_subtile_3__pin_sc_in_0_),
		.left_width_0_height_0_subtile_3__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_3__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_3__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_3__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_3__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_3__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_4__pin_f2a_i_0_(cby_9__1__0_right_grid_left_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_4__pin_sc_in_0_(grid_io_right_10__1__undriven_left_width_0_height_0_subtile_4__pin_sc_in_0_),
		.left_width_0_height_0_subtile_4__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_4__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_4__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_4__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_4__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_4__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_5__pin_f2a_i_0_(cby_9__1__0_right_grid_left_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_5__pin_sc_in_0_(grid_io_right_10__1__undriven_left_width_0_height_0_subtile_5__pin_sc_in_0_),
		.left_width_0_height_0_subtile_5__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_5__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_5__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_5__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_5__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_5__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_6__pin_f2a_i_0_(cby_9__1__0_right_grid_left_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_6__pin_sc_in_0_(grid_io_right_10__1__undriven_left_width_0_height_0_subtile_6__pin_sc_in_0_),
		.left_width_0_height_0_subtile_6__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_6__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_6__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_6__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_6__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_6__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_7__pin_f2a_i_0_(cby_9__1__0_right_grid_left_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_7__pin_sc_in_0_(grid_io_right_10__1__undriven_left_width_0_height_0_subtile_7__pin_sc_in_0_),
		.left_width_0_height_0_subtile_7__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_7__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_7__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_7__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_7__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_7__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_8__pin_f2a_i_0_(cby_9__1__0_right_grid_left_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_8__pin_sc_in_0_(grid_io_right_10__1__undriven_left_width_0_height_0_subtile_8__pin_sc_in_0_),
		.left_width_0_height_0_subtile_8__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_8__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_8__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_8__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_8__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_8__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_9__pin_f2a_i_0_(cby_9__1__0_right_grid_left_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_9__pin_sc_in_0_(grid_io_right_10__1__undriven_left_width_0_height_0_subtile_9__pin_sc_in_0_),
		.left_width_0_height_0_subtile_9__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_9__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_9__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_9__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_9__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_9__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_10__pin_f2a_i_0_(cby_9__1__0_right_grid_left_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_10__pin_sc_in_0_(grid_io_right_10__1__undriven_left_width_0_height_0_subtile_10__pin_sc_in_0_),
		.left_width_0_height_0_subtile_10__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_10__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_10__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_10__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_10__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_10__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_11__pin_f2a_i_0_(cby_9__1__0_right_grid_left_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_11__pin_sc_in_0_(grid_io_right_10__1__undriven_left_width_0_height_0_subtile_11__pin_sc_in_0_),
		.left_width_0_height_0_subtile_11__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_11__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_11__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_11__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_11__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_11__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_12__pin_f2a_i_0_(cby_9__1__0_right_grid_left_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_12__pin_sc_in_0_(grid_io_right_10__1__undriven_left_width_0_height_0_subtile_12__pin_sc_in_0_),
		.left_width_0_height_0_subtile_12__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_12__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_12__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_12__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_12__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_12__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_13__pin_f2a_i_0_(cby_9__1__0_right_grid_left_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_13__pin_sc_in_0_(grid_io_right_10__1__undriven_left_width_0_height_0_subtile_13__pin_sc_in_0_),
		.left_width_0_height_0_subtile_13__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_13__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_13__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_13__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_13__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_13__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_14__pin_f2a_i_0_(cby_9__1__0_right_grid_left_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_14__pin_sc_in_0_(grid_io_right_10__1__undriven_left_width_0_height_0_subtile_14__pin_sc_in_0_),
		.left_width_0_height_0_subtile_14__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_14__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_14__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_14__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_14__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_14__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_15__pin_f2a_i_0_(cby_9__1__0_right_grid_left_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_15__pin_sc_in_0_(grid_io_right_10__1__undriven_left_width_0_height_0_subtile_15__pin_sc_in_0_),
		.left_width_0_height_0_subtile_15__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_15__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_15__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_15__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_15__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_15__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_16__pin_f2a_i_0_(cby_9__1__0_right_grid_left_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_16__pin_sc_in_0_(grid_io_right_10__1__undriven_left_width_0_height_0_subtile_16__pin_sc_in_0_),
		.left_width_0_height_0_subtile_16__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_16__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_16__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_16__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_16__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_16__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_17__pin_f2a_i_0_(cby_9__1__0_right_grid_left_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_17__pin_sc_in_0_(grid_io_right_10__1__undriven_left_width_0_height_0_subtile_17__pin_sc_in_0_),
		.left_width_0_height_0_subtile_17__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_17__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_17__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_17__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_17__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_17__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_18__pin_f2a_i_0_(cby_9__1__0_right_grid_left_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_18__pin_sc_in_0_(grid_io_right_10__1__undriven_left_width_0_height_0_subtile_18__pin_sc_in_0_),
		.left_width_0_height_0_subtile_18__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_18__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_18__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_18__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_18__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_18__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_19__pin_f2a_i_0_(cby_9__1__0_right_grid_left_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_19__pin_sc_in_0_(grid_io_right_10__1__undriven_left_width_0_height_0_subtile_19__pin_sc_in_0_),
		.left_width_0_height_0_subtile_19__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_19__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_19__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_19__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_19__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_19__pin_clk_3_(clk[3]),
		.ccff_head(grid_io_bottom_7_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_0__pin_sc_out_0_(grid_io_right_10__1__undriven_left_width_0_height_0_subtile_0__pin_sc_out_0_),
		.left_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_1__pin_sc_out_0_(grid_io_right_10__1__undriven_left_width_0_height_0_subtile_1__pin_sc_out_0_),
		.left_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_2__pin_sc_out_0_(grid_io_right_10__1__undriven_left_width_0_height_0_subtile_2__pin_sc_out_0_),
		.left_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_3__pin_sc_out_0_(grid_io_right_10__1__undriven_left_width_0_height_0_subtile_3__pin_sc_out_0_),
		.left_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_4__pin_sc_out_0_(grid_io_right_10__1__undriven_left_width_0_height_0_subtile_4__pin_sc_out_0_),
		.left_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_5__pin_sc_out_0_(grid_io_right_10__1__undriven_left_width_0_height_0_subtile_5__pin_sc_out_0_),
		.left_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_6__pin_sc_out_0_(grid_io_right_10__1__undriven_left_width_0_height_0_subtile_6__pin_sc_out_0_),
		.left_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_7__pin_sc_out_0_(grid_io_right_10__1__undriven_left_width_0_height_0_subtile_7__pin_sc_out_0_),
		.left_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_8__pin_sc_out_0_(grid_io_right_10__1__undriven_left_width_0_height_0_subtile_8__pin_sc_out_0_),
		.left_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_9__pin_sc_out_0_(grid_io_right_10__1__undriven_left_width_0_height_0_subtile_9__pin_sc_out_0_),
		.left_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_10__pin_sc_out_0_(grid_io_right_10__1__undriven_left_width_0_height_0_subtile_10__pin_sc_out_0_),
		.left_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_11__pin_sc_out_0_(grid_io_right_10__1__undriven_left_width_0_height_0_subtile_11__pin_sc_out_0_),
		.left_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_12__pin_sc_out_0_(grid_io_right_10__1__undriven_left_width_0_height_0_subtile_12__pin_sc_out_0_),
		.left_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_13__pin_sc_out_0_(grid_io_right_10__1__undriven_left_width_0_height_0_subtile_13__pin_sc_out_0_),
		.left_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_14__pin_sc_out_0_(grid_io_right_10__1__undriven_left_width_0_height_0_subtile_14__pin_sc_out_0_),
		.left_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_15__pin_sc_out_0_(grid_io_right_10__1__undriven_left_width_0_height_0_subtile_15__pin_sc_out_0_),
		.left_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_16__pin_sc_out_0_(grid_io_right_10__1__undriven_left_width_0_height_0_subtile_16__pin_sc_out_0_),
		.left_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_17__pin_sc_out_0_(grid_io_right_10__1__undriven_left_width_0_height_0_subtile_17__pin_sc_out_0_),
		.left_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_18__pin_sc_out_0_(grid_io_right_10__1__undriven_left_width_0_height_0_subtile_18__pin_sc_out_0_),
		.left_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_19__pin_sc_out_0_(grid_io_right_10__1__undriven_left_width_0_height_0_subtile_19__pin_sc_out_0_),
		.ccff_tail(grid_io_right_0_ccff_tail));

	grid_io_right grid_io_right_10__2_ (
		.test_en(test_en),
		.scan_mode(scan_mode),
		.scan_clk(scan_clk),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.CFG_DONE(CFG_DONE),
		.gfpga_pad_QL_PREIO_A2F(gfpga_pad_QL_PREIO_A2F[440:459]),
		.gfpga_pad_QL_PREIO_F2A(gfpga_pad_QL_PREIO_F2A[440:459]),
		.gfpga_pad_QL_PREIO_F2A_DEF0(gfpga_pad_QL_PREIO_F2A_DEF0[440:459]),
		.gfpga_pad_QL_PREIO_F2A_DEF1(gfpga_pad_QL_PREIO_F2A_DEF1[440:459]),
		.gfpga_pad_QL_PREIO_F2A_CLK(gfpga_pad_QL_PREIO_F2A_CLK[440:459]),
		.left_width_0_height_0_subtile_0__pin_f2a_i_0_(cby_9__2__0_right_grid_left_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_0__pin_sc_in_0_(grid_io_right_10__2__undriven_left_width_0_height_0_subtile_0__pin_sc_in_0_),
		.left_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_1__pin_f2a_i_0_(cby_9__2__0_right_grid_left_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_1__pin_sc_in_0_(grid_io_right_10__2__undriven_left_width_0_height_0_subtile_1__pin_sc_in_0_),
		.left_width_0_height_0_subtile_1__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_1__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_1__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_1__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_1__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_1__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_2__pin_f2a_i_0_(cby_9__2__0_right_grid_left_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_2__pin_sc_in_0_(grid_io_right_10__2__undriven_left_width_0_height_0_subtile_2__pin_sc_in_0_),
		.left_width_0_height_0_subtile_2__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_2__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_2__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_2__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_2__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_2__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_3__pin_f2a_i_0_(cby_9__2__0_right_grid_left_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_3__pin_sc_in_0_(grid_io_right_10__2__undriven_left_width_0_height_0_subtile_3__pin_sc_in_0_),
		.left_width_0_height_0_subtile_3__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_3__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_3__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_3__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_3__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_3__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_4__pin_f2a_i_0_(cby_9__2__0_right_grid_left_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_4__pin_sc_in_0_(grid_io_right_10__2__undriven_left_width_0_height_0_subtile_4__pin_sc_in_0_),
		.left_width_0_height_0_subtile_4__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_4__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_4__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_4__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_4__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_4__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_5__pin_f2a_i_0_(cby_9__2__0_right_grid_left_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_5__pin_sc_in_0_(grid_io_right_10__2__undriven_left_width_0_height_0_subtile_5__pin_sc_in_0_),
		.left_width_0_height_0_subtile_5__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_5__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_5__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_5__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_5__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_5__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_6__pin_f2a_i_0_(cby_9__2__0_right_grid_left_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_6__pin_sc_in_0_(grid_io_right_10__2__undriven_left_width_0_height_0_subtile_6__pin_sc_in_0_),
		.left_width_0_height_0_subtile_6__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_6__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_6__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_6__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_6__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_6__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_7__pin_f2a_i_0_(cby_9__2__0_right_grid_left_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_7__pin_sc_in_0_(grid_io_right_10__2__undriven_left_width_0_height_0_subtile_7__pin_sc_in_0_),
		.left_width_0_height_0_subtile_7__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_7__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_7__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_7__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_7__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_7__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_8__pin_f2a_i_0_(cby_9__2__0_right_grid_left_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_8__pin_sc_in_0_(grid_io_right_10__2__undriven_left_width_0_height_0_subtile_8__pin_sc_in_0_),
		.left_width_0_height_0_subtile_8__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_8__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_8__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_8__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_8__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_8__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_9__pin_f2a_i_0_(cby_9__2__0_right_grid_left_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_9__pin_sc_in_0_(grid_io_right_10__2__undriven_left_width_0_height_0_subtile_9__pin_sc_in_0_),
		.left_width_0_height_0_subtile_9__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_9__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_9__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_9__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_9__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_9__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_10__pin_f2a_i_0_(cby_9__2__0_right_grid_left_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_10__pin_sc_in_0_(grid_io_right_10__2__undriven_left_width_0_height_0_subtile_10__pin_sc_in_0_),
		.left_width_0_height_0_subtile_10__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_10__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_10__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_10__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_10__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_10__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_11__pin_f2a_i_0_(cby_9__2__0_right_grid_left_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_11__pin_sc_in_0_(grid_io_right_10__2__undriven_left_width_0_height_0_subtile_11__pin_sc_in_0_),
		.left_width_0_height_0_subtile_11__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_11__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_11__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_11__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_11__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_11__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_12__pin_f2a_i_0_(cby_9__2__0_right_grid_left_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_12__pin_sc_in_0_(grid_io_right_10__2__undriven_left_width_0_height_0_subtile_12__pin_sc_in_0_),
		.left_width_0_height_0_subtile_12__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_12__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_12__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_12__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_12__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_12__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_13__pin_f2a_i_0_(cby_9__2__0_right_grid_left_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_13__pin_sc_in_0_(grid_io_right_10__2__undriven_left_width_0_height_0_subtile_13__pin_sc_in_0_),
		.left_width_0_height_0_subtile_13__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_13__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_13__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_13__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_13__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_13__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_14__pin_f2a_i_0_(cby_9__2__0_right_grid_left_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_14__pin_sc_in_0_(grid_io_right_10__2__undriven_left_width_0_height_0_subtile_14__pin_sc_in_0_),
		.left_width_0_height_0_subtile_14__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_14__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_14__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_14__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_14__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_14__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_15__pin_f2a_i_0_(cby_9__2__0_right_grid_left_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_15__pin_sc_in_0_(grid_io_right_10__2__undriven_left_width_0_height_0_subtile_15__pin_sc_in_0_),
		.left_width_0_height_0_subtile_15__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_15__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_15__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_15__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_15__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_15__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_16__pin_f2a_i_0_(cby_9__2__0_right_grid_left_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_16__pin_sc_in_0_(grid_io_right_10__2__undriven_left_width_0_height_0_subtile_16__pin_sc_in_0_),
		.left_width_0_height_0_subtile_16__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_16__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_16__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_16__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_16__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_16__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_17__pin_f2a_i_0_(cby_9__2__0_right_grid_left_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_17__pin_sc_in_0_(grid_io_right_10__2__undriven_left_width_0_height_0_subtile_17__pin_sc_in_0_),
		.left_width_0_height_0_subtile_17__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_17__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_17__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_17__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_17__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_17__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_18__pin_f2a_i_0_(cby_9__2__0_right_grid_left_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_18__pin_sc_in_0_(grid_io_right_10__2__undriven_left_width_0_height_0_subtile_18__pin_sc_in_0_),
		.left_width_0_height_0_subtile_18__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_18__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_18__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_18__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_18__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_18__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_19__pin_f2a_i_0_(cby_9__2__0_right_grid_left_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_19__pin_sc_in_0_(grid_io_right_10__2__undriven_left_width_0_height_0_subtile_19__pin_sc_in_0_),
		.left_width_0_height_0_subtile_19__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_19__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_19__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_19__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_19__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_19__pin_clk_3_(clk[3]),
		.ccff_head(sb_10__1__0_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_0__pin_sc_out_0_(grid_io_right_10__2__undriven_left_width_0_height_0_subtile_0__pin_sc_out_0_),
		.left_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_1__pin_sc_out_0_(grid_io_right_10__2__undriven_left_width_0_height_0_subtile_1__pin_sc_out_0_),
		.left_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_2__pin_sc_out_0_(grid_io_right_10__2__undriven_left_width_0_height_0_subtile_2__pin_sc_out_0_),
		.left_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_3__pin_sc_out_0_(grid_io_right_10__2__undriven_left_width_0_height_0_subtile_3__pin_sc_out_0_),
		.left_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_4__pin_sc_out_0_(grid_io_right_10__2__undriven_left_width_0_height_0_subtile_4__pin_sc_out_0_),
		.left_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_5__pin_sc_out_0_(grid_io_right_10__2__undriven_left_width_0_height_0_subtile_5__pin_sc_out_0_),
		.left_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_6__pin_sc_out_0_(grid_io_right_10__2__undriven_left_width_0_height_0_subtile_6__pin_sc_out_0_),
		.left_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_7__pin_sc_out_0_(grid_io_right_10__2__undriven_left_width_0_height_0_subtile_7__pin_sc_out_0_),
		.left_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_8__pin_sc_out_0_(grid_io_right_10__2__undriven_left_width_0_height_0_subtile_8__pin_sc_out_0_),
		.left_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_9__pin_sc_out_0_(grid_io_right_10__2__undriven_left_width_0_height_0_subtile_9__pin_sc_out_0_),
		.left_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_10__pin_sc_out_0_(grid_io_right_10__2__undriven_left_width_0_height_0_subtile_10__pin_sc_out_0_),
		.left_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_11__pin_sc_out_0_(grid_io_right_10__2__undriven_left_width_0_height_0_subtile_11__pin_sc_out_0_),
		.left_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_12__pin_sc_out_0_(grid_io_right_10__2__undriven_left_width_0_height_0_subtile_12__pin_sc_out_0_),
		.left_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_13__pin_sc_out_0_(grid_io_right_10__2__undriven_left_width_0_height_0_subtile_13__pin_sc_out_0_),
		.left_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_14__pin_sc_out_0_(grid_io_right_10__2__undriven_left_width_0_height_0_subtile_14__pin_sc_out_0_),
		.left_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_15__pin_sc_out_0_(grid_io_right_10__2__undriven_left_width_0_height_0_subtile_15__pin_sc_out_0_),
		.left_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_16__pin_sc_out_0_(grid_io_right_10__2__undriven_left_width_0_height_0_subtile_16__pin_sc_out_0_),
		.left_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_17__pin_sc_out_0_(grid_io_right_10__2__undriven_left_width_0_height_0_subtile_17__pin_sc_out_0_),
		.left_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_18__pin_sc_out_0_(grid_io_right_10__2__undriven_left_width_0_height_0_subtile_18__pin_sc_out_0_),
		.left_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_19__pin_sc_out_0_(grid_io_right_10__2__undriven_left_width_0_height_0_subtile_19__pin_sc_out_0_),
		.ccff_tail(grid_io_right_1_ccff_tail));

	grid_io_right grid_io_right_10__3_ (
		.test_en(test_en),
		.scan_mode(scan_mode),
		.scan_clk(scan_clk),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.CFG_DONE(CFG_DONE),
		.gfpga_pad_QL_PREIO_A2F(gfpga_pad_QL_PREIO_A2F[420:439]),
		.gfpga_pad_QL_PREIO_F2A(gfpga_pad_QL_PREIO_F2A[420:439]),
		.gfpga_pad_QL_PREIO_F2A_DEF0(gfpga_pad_QL_PREIO_F2A_DEF0[420:439]),
		.gfpga_pad_QL_PREIO_F2A_DEF1(gfpga_pad_QL_PREIO_F2A_DEF1[420:439]),
		.gfpga_pad_QL_PREIO_F2A_CLK(gfpga_pad_QL_PREIO_F2A_CLK[420:439]),
		.left_width_0_height_0_subtile_0__pin_f2a_i_0_(cby_9__2__1_right_grid_left_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_0__pin_sc_in_0_(grid_io_right_10__3__undriven_left_width_0_height_0_subtile_0__pin_sc_in_0_),
		.left_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_1__pin_f2a_i_0_(cby_9__2__1_right_grid_left_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_1__pin_sc_in_0_(grid_io_right_10__3__undriven_left_width_0_height_0_subtile_1__pin_sc_in_0_),
		.left_width_0_height_0_subtile_1__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_1__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_1__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_1__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_1__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_1__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_2__pin_f2a_i_0_(cby_9__2__1_right_grid_left_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_2__pin_sc_in_0_(grid_io_right_10__3__undriven_left_width_0_height_0_subtile_2__pin_sc_in_0_),
		.left_width_0_height_0_subtile_2__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_2__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_2__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_2__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_2__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_2__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_3__pin_f2a_i_0_(cby_9__2__1_right_grid_left_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_3__pin_sc_in_0_(grid_io_right_10__3__undriven_left_width_0_height_0_subtile_3__pin_sc_in_0_),
		.left_width_0_height_0_subtile_3__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_3__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_3__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_3__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_3__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_3__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_4__pin_f2a_i_0_(cby_9__2__1_right_grid_left_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_4__pin_sc_in_0_(grid_io_right_10__3__undriven_left_width_0_height_0_subtile_4__pin_sc_in_0_),
		.left_width_0_height_0_subtile_4__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_4__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_4__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_4__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_4__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_4__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_5__pin_f2a_i_0_(cby_9__2__1_right_grid_left_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_5__pin_sc_in_0_(grid_io_right_10__3__undriven_left_width_0_height_0_subtile_5__pin_sc_in_0_),
		.left_width_0_height_0_subtile_5__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_5__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_5__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_5__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_5__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_5__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_6__pin_f2a_i_0_(cby_9__2__1_right_grid_left_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_6__pin_sc_in_0_(grid_io_right_10__3__undriven_left_width_0_height_0_subtile_6__pin_sc_in_0_),
		.left_width_0_height_0_subtile_6__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_6__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_6__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_6__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_6__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_6__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_7__pin_f2a_i_0_(cby_9__2__1_right_grid_left_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_7__pin_sc_in_0_(grid_io_right_10__3__undriven_left_width_0_height_0_subtile_7__pin_sc_in_0_),
		.left_width_0_height_0_subtile_7__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_7__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_7__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_7__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_7__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_7__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_8__pin_f2a_i_0_(cby_9__2__1_right_grid_left_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_8__pin_sc_in_0_(grid_io_right_10__3__undriven_left_width_0_height_0_subtile_8__pin_sc_in_0_),
		.left_width_0_height_0_subtile_8__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_8__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_8__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_8__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_8__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_8__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_9__pin_f2a_i_0_(cby_9__2__1_right_grid_left_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_9__pin_sc_in_0_(grid_io_right_10__3__undriven_left_width_0_height_0_subtile_9__pin_sc_in_0_),
		.left_width_0_height_0_subtile_9__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_9__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_9__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_9__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_9__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_9__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_10__pin_f2a_i_0_(cby_9__2__1_right_grid_left_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_10__pin_sc_in_0_(grid_io_right_10__3__undriven_left_width_0_height_0_subtile_10__pin_sc_in_0_),
		.left_width_0_height_0_subtile_10__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_10__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_10__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_10__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_10__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_10__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_11__pin_f2a_i_0_(cby_9__2__1_right_grid_left_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_11__pin_sc_in_0_(grid_io_right_10__3__undriven_left_width_0_height_0_subtile_11__pin_sc_in_0_),
		.left_width_0_height_0_subtile_11__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_11__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_11__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_11__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_11__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_11__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_12__pin_f2a_i_0_(cby_9__2__1_right_grid_left_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_12__pin_sc_in_0_(grid_io_right_10__3__undriven_left_width_0_height_0_subtile_12__pin_sc_in_0_),
		.left_width_0_height_0_subtile_12__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_12__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_12__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_12__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_12__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_12__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_13__pin_f2a_i_0_(cby_9__2__1_right_grid_left_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_13__pin_sc_in_0_(grid_io_right_10__3__undriven_left_width_0_height_0_subtile_13__pin_sc_in_0_),
		.left_width_0_height_0_subtile_13__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_13__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_13__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_13__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_13__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_13__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_14__pin_f2a_i_0_(cby_9__2__1_right_grid_left_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_14__pin_sc_in_0_(grid_io_right_10__3__undriven_left_width_0_height_0_subtile_14__pin_sc_in_0_),
		.left_width_0_height_0_subtile_14__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_14__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_14__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_14__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_14__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_14__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_15__pin_f2a_i_0_(cby_9__2__1_right_grid_left_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_15__pin_sc_in_0_(grid_io_right_10__3__undriven_left_width_0_height_0_subtile_15__pin_sc_in_0_),
		.left_width_0_height_0_subtile_15__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_15__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_15__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_15__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_15__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_15__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_16__pin_f2a_i_0_(cby_9__2__1_right_grid_left_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_16__pin_sc_in_0_(grid_io_right_10__3__undriven_left_width_0_height_0_subtile_16__pin_sc_in_0_),
		.left_width_0_height_0_subtile_16__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_16__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_16__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_16__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_16__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_16__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_17__pin_f2a_i_0_(cby_9__2__1_right_grid_left_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_17__pin_sc_in_0_(grid_io_right_10__3__undriven_left_width_0_height_0_subtile_17__pin_sc_in_0_),
		.left_width_0_height_0_subtile_17__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_17__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_17__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_17__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_17__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_17__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_18__pin_f2a_i_0_(cby_9__2__1_right_grid_left_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_18__pin_sc_in_0_(grid_io_right_10__3__undriven_left_width_0_height_0_subtile_18__pin_sc_in_0_),
		.left_width_0_height_0_subtile_18__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_18__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_18__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_18__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_18__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_18__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_19__pin_f2a_i_0_(cby_9__2__1_right_grid_left_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_19__pin_sc_in_0_(grid_io_right_10__3__undriven_left_width_0_height_0_subtile_19__pin_sc_in_0_),
		.left_width_0_height_0_subtile_19__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_19__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_19__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_19__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_19__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_19__pin_clk_3_(clk[3]),
		.ccff_head(sb_10__1__1_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_0__pin_sc_out_0_(grid_io_right_10__3__undriven_left_width_0_height_0_subtile_0__pin_sc_out_0_),
		.left_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_1__pin_sc_out_0_(grid_io_right_10__3__undriven_left_width_0_height_0_subtile_1__pin_sc_out_0_),
		.left_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_2__pin_sc_out_0_(grid_io_right_10__3__undriven_left_width_0_height_0_subtile_2__pin_sc_out_0_),
		.left_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_3__pin_sc_out_0_(grid_io_right_10__3__undriven_left_width_0_height_0_subtile_3__pin_sc_out_0_),
		.left_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_4__pin_sc_out_0_(grid_io_right_10__3__undriven_left_width_0_height_0_subtile_4__pin_sc_out_0_),
		.left_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_5__pin_sc_out_0_(grid_io_right_10__3__undriven_left_width_0_height_0_subtile_5__pin_sc_out_0_),
		.left_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_6__pin_sc_out_0_(grid_io_right_10__3__undriven_left_width_0_height_0_subtile_6__pin_sc_out_0_),
		.left_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_7__pin_sc_out_0_(grid_io_right_10__3__undriven_left_width_0_height_0_subtile_7__pin_sc_out_0_),
		.left_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_8__pin_sc_out_0_(grid_io_right_10__3__undriven_left_width_0_height_0_subtile_8__pin_sc_out_0_),
		.left_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_9__pin_sc_out_0_(grid_io_right_10__3__undriven_left_width_0_height_0_subtile_9__pin_sc_out_0_),
		.left_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_10__pin_sc_out_0_(grid_io_right_10__3__undriven_left_width_0_height_0_subtile_10__pin_sc_out_0_),
		.left_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_11__pin_sc_out_0_(grid_io_right_10__3__undriven_left_width_0_height_0_subtile_11__pin_sc_out_0_),
		.left_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_12__pin_sc_out_0_(grid_io_right_10__3__undriven_left_width_0_height_0_subtile_12__pin_sc_out_0_),
		.left_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_13__pin_sc_out_0_(grid_io_right_10__3__undriven_left_width_0_height_0_subtile_13__pin_sc_out_0_),
		.left_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_14__pin_sc_out_0_(grid_io_right_10__3__undriven_left_width_0_height_0_subtile_14__pin_sc_out_0_),
		.left_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_15__pin_sc_out_0_(grid_io_right_10__3__undriven_left_width_0_height_0_subtile_15__pin_sc_out_0_),
		.left_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_16__pin_sc_out_0_(grid_io_right_10__3__undriven_left_width_0_height_0_subtile_16__pin_sc_out_0_),
		.left_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_17__pin_sc_out_0_(grid_io_right_10__3__undriven_left_width_0_height_0_subtile_17__pin_sc_out_0_),
		.left_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_18__pin_sc_out_0_(grid_io_right_10__3__undriven_left_width_0_height_0_subtile_18__pin_sc_out_0_),
		.left_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_19__pin_sc_out_0_(grid_io_right_10__3__undriven_left_width_0_height_0_subtile_19__pin_sc_out_0_),
		.ccff_tail(grid_io_right_2_ccff_tail));

	grid_io_right grid_io_right_10__4_ (
		.test_en(test_en),
		.scan_mode(scan_mode),
		.scan_clk(scan_clk),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.CFG_DONE(CFG_DONE),
		.gfpga_pad_QL_PREIO_A2F(gfpga_pad_QL_PREIO_A2F[400:419]),
		.gfpga_pad_QL_PREIO_F2A(gfpga_pad_QL_PREIO_F2A[400:419]),
		.gfpga_pad_QL_PREIO_F2A_DEF0(gfpga_pad_QL_PREIO_F2A_DEF0[400:419]),
		.gfpga_pad_QL_PREIO_F2A_DEF1(gfpga_pad_QL_PREIO_F2A_DEF1[400:419]),
		.gfpga_pad_QL_PREIO_F2A_CLK(gfpga_pad_QL_PREIO_F2A_CLK[400:419]),
		.left_width_0_height_0_subtile_0__pin_f2a_i_0_(cby_9__2__2_right_grid_left_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_0__pin_sc_in_0_(grid_io_right_10__4__undriven_left_width_0_height_0_subtile_0__pin_sc_in_0_),
		.left_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_1__pin_f2a_i_0_(cby_9__2__2_right_grid_left_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_1__pin_sc_in_0_(grid_io_right_10__4__undriven_left_width_0_height_0_subtile_1__pin_sc_in_0_),
		.left_width_0_height_0_subtile_1__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_1__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_1__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_1__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_1__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_1__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_2__pin_f2a_i_0_(cby_9__2__2_right_grid_left_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_2__pin_sc_in_0_(grid_io_right_10__4__undriven_left_width_0_height_0_subtile_2__pin_sc_in_0_),
		.left_width_0_height_0_subtile_2__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_2__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_2__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_2__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_2__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_2__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_3__pin_f2a_i_0_(cby_9__2__2_right_grid_left_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_3__pin_sc_in_0_(grid_io_right_10__4__undriven_left_width_0_height_0_subtile_3__pin_sc_in_0_),
		.left_width_0_height_0_subtile_3__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_3__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_3__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_3__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_3__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_3__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_4__pin_f2a_i_0_(cby_9__2__2_right_grid_left_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_4__pin_sc_in_0_(grid_io_right_10__4__undriven_left_width_0_height_0_subtile_4__pin_sc_in_0_),
		.left_width_0_height_0_subtile_4__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_4__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_4__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_4__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_4__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_4__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_5__pin_f2a_i_0_(cby_9__2__2_right_grid_left_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_5__pin_sc_in_0_(grid_io_right_10__4__undriven_left_width_0_height_0_subtile_5__pin_sc_in_0_),
		.left_width_0_height_0_subtile_5__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_5__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_5__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_5__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_5__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_5__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_6__pin_f2a_i_0_(cby_9__2__2_right_grid_left_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_6__pin_sc_in_0_(grid_io_right_10__4__undriven_left_width_0_height_0_subtile_6__pin_sc_in_0_),
		.left_width_0_height_0_subtile_6__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_6__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_6__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_6__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_6__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_6__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_7__pin_f2a_i_0_(cby_9__2__2_right_grid_left_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_7__pin_sc_in_0_(grid_io_right_10__4__undriven_left_width_0_height_0_subtile_7__pin_sc_in_0_),
		.left_width_0_height_0_subtile_7__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_7__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_7__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_7__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_7__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_7__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_8__pin_f2a_i_0_(cby_9__2__2_right_grid_left_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_8__pin_sc_in_0_(grid_io_right_10__4__undriven_left_width_0_height_0_subtile_8__pin_sc_in_0_),
		.left_width_0_height_0_subtile_8__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_8__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_8__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_8__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_8__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_8__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_9__pin_f2a_i_0_(cby_9__2__2_right_grid_left_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_9__pin_sc_in_0_(grid_io_right_10__4__undriven_left_width_0_height_0_subtile_9__pin_sc_in_0_),
		.left_width_0_height_0_subtile_9__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_9__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_9__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_9__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_9__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_9__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_10__pin_f2a_i_0_(cby_9__2__2_right_grid_left_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_10__pin_sc_in_0_(grid_io_right_10__4__undriven_left_width_0_height_0_subtile_10__pin_sc_in_0_),
		.left_width_0_height_0_subtile_10__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_10__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_10__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_10__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_10__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_10__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_11__pin_f2a_i_0_(cby_9__2__2_right_grid_left_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_11__pin_sc_in_0_(grid_io_right_10__4__undriven_left_width_0_height_0_subtile_11__pin_sc_in_0_),
		.left_width_0_height_0_subtile_11__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_11__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_11__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_11__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_11__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_11__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_12__pin_f2a_i_0_(cby_9__2__2_right_grid_left_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_12__pin_sc_in_0_(grid_io_right_10__4__undriven_left_width_0_height_0_subtile_12__pin_sc_in_0_),
		.left_width_0_height_0_subtile_12__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_12__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_12__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_12__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_12__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_12__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_13__pin_f2a_i_0_(cby_9__2__2_right_grid_left_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_13__pin_sc_in_0_(grid_io_right_10__4__undriven_left_width_0_height_0_subtile_13__pin_sc_in_0_),
		.left_width_0_height_0_subtile_13__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_13__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_13__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_13__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_13__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_13__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_14__pin_f2a_i_0_(cby_9__2__2_right_grid_left_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_14__pin_sc_in_0_(grid_io_right_10__4__undriven_left_width_0_height_0_subtile_14__pin_sc_in_0_),
		.left_width_0_height_0_subtile_14__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_14__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_14__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_14__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_14__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_14__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_15__pin_f2a_i_0_(cby_9__2__2_right_grid_left_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_15__pin_sc_in_0_(grid_io_right_10__4__undriven_left_width_0_height_0_subtile_15__pin_sc_in_0_),
		.left_width_0_height_0_subtile_15__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_15__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_15__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_15__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_15__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_15__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_16__pin_f2a_i_0_(cby_9__2__2_right_grid_left_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_16__pin_sc_in_0_(grid_io_right_10__4__undriven_left_width_0_height_0_subtile_16__pin_sc_in_0_),
		.left_width_0_height_0_subtile_16__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_16__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_16__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_16__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_16__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_16__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_17__pin_f2a_i_0_(cby_9__2__2_right_grid_left_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_17__pin_sc_in_0_(grid_io_right_10__4__undriven_left_width_0_height_0_subtile_17__pin_sc_in_0_),
		.left_width_0_height_0_subtile_17__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_17__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_17__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_17__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_17__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_17__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_18__pin_f2a_i_0_(cby_9__2__2_right_grid_left_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_18__pin_sc_in_0_(grid_io_right_10__4__undriven_left_width_0_height_0_subtile_18__pin_sc_in_0_),
		.left_width_0_height_0_subtile_18__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_18__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_18__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_18__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_18__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_18__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_19__pin_f2a_i_0_(cby_9__2__2_right_grid_left_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_19__pin_sc_in_0_(grid_io_right_10__4__undriven_left_width_0_height_0_subtile_19__pin_sc_in_0_),
		.left_width_0_height_0_subtile_19__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_19__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_19__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_19__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_19__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_19__pin_clk_3_(clk[3]),
		.ccff_head(ccff_head[4]),
		.left_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_0__pin_sc_out_0_(grid_io_right_10__4__undriven_left_width_0_height_0_subtile_0__pin_sc_out_0_),
		.left_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_1__pin_sc_out_0_(grid_io_right_10__4__undriven_left_width_0_height_0_subtile_1__pin_sc_out_0_),
		.left_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_2__pin_sc_out_0_(grid_io_right_10__4__undriven_left_width_0_height_0_subtile_2__pin_sc_out_0_),
		.left_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_3__pin_sc_out_0_(grid_io_right_10__4__undriven_left_width_0_height_0_subtile_3__pin_sc_out_0_),
		.left_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_4__pin_sc_out_0_(grid_io_right_10__4__undriven_left_width_0_height_0_subtile_4__pin_sc_out_0_),
		.left_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_5__pin_sc_out_0_(grid_io_right_10__4__undriven_left_width_0_height_0_subtile_5__pin_sc_out_0_),
		.left_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_6__pin_sc_out_0_(grid_io_right_10__4__undriven_left_width_0_height_0_subtile_6__pin_sc_out_0_),
		.left_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_7__pin_sc_out_0_(grid_io_right_10__4__undriven_left_width_0_height_0_subtile_7__pin_sc_out_0_),
		.left_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_8__pin_sc_out_0_(grid_io_right_10__4__undriven_left_width_0_height_0_subtile_8__pin_sc_out_0_),
		.left_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_9__pin_sc_out_0_(grid_io_right_10__4__undriven_left_width_0_height_0_subtile_9__pin_sc_out_0_),
		.left_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_10__pin_sc_out_0_(grid_io_right_10__4__undriven_left_width_0_height_0_subtile_10__pin_sc_out_0_),
		.left_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_11__pin_sc_out_0_(grid_io_right_10__4__undriven_left_width_0_height_0_subtile_11__pin_sc_out_0_),
		.left_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_12__pin_sc_out_0_(grid_io_right_10__4__undriven_left_width_0_height_0_subtile_12__pin_sc_out_0_),
		.left_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_13__pin_sc_out_0_(grid_io_right_10__4__undriven_left_width_0_height_0_subtile_13__pin_sc_out_0_),
		.left_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_14__pin_sc_out_0_(grid_io_right_10__4__undriven_left_width_0_height_0_subtile_14__pin_sc_out_0_),
		.left_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_15__pin_sc_out_0_(grid_io_right_10__4__undriven_left_width_0_height_0_subtile_15__pin_sc_out_0_),
		.left_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_16__pin_sc_out_0_(grid_io_right_10__4__undriven_left_width_0_height_0_subtile_16__pin_sc_out_0_),
		.left_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_17__pin_sc_out_0_(grid_io_right_10__4__undriven_left_width_0_height_0_subtile_17__pin_sc_out_0_),
		.left_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_18__pin_sc_out_0_(grid_io_right_10__4__undriven_left_width_0_height_0_subtile_18__pin_sc_out_0_),
		.left_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_19__pin_sc_out_0_(grid_io_right_10__4__undriven_left_width_0_height_0_subtile_19__pin_sc_out_0_),
		.ccff_tail(grid_io_right_3_ccff_tail));

	grid_io_right grid_io_right_10__5_ (
		.test_en(test_en),
		.scan_mode(scan_mode),
		.scan_clk(scan_clk),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.CFG_DONE(CFG_DONE),
		.gfpga_pad_QL_PREIO_A2F(gfpga_pad_QL_PREIO_A2F[380:399]),
		.gfpga_pad_QL_PREIO_F2A(gfpga_pad_QL_PREIO_F2A[380:399]),
		.gfpga_pad_QL_PREIO_F2A_DEF0(gfpga_pad_QL_PREIO_F2A_DEF0[380:399]),
		.gfpga_pad_QL_PREIO_F2A_DEF1(gfpga_pad_QL_PREIO_F2A_DEF1[380:399]),
		.gfpga_pad_QL_PREIO_F2A_CLK(gfpga_pad_QL_PREIO_F2A_CLK[380:399]),
		.left_width_0_height_0_subtile_0__pin_f2a_i_0_(cby_9__2__3_right_grid_left_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_0__pin_sc_in_0_(grid_io_right_10__5__undriven_left_width_0_height_0_subtile_0__pin_sc_in_0_),
		.left_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_1__pin_f2a_i_0_(cby_9__2__3_right_grid_left_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_1__pin_sc_in_0_(grid_io_right_10__5__undriven_left_width_0_height_0_subtile_1__pin_sc_in_0_),
		.left_width_0_height_0_subtile_1__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_1__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_1__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_1__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_1__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_1__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_2__pin_f2a_i_0_(cby_9__2__3_right_grid_left_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_2__pin_sc_in_0_(grid_io_right_10__5__undriven_left_width_0_height_0_subtile_2__pin_sc_in_0_),
		.left_width_0_height_0_subtile_2__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_2__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_2__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_2__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_2__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_2__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_3__pin_f2a_i_0_(cby_9__2__3_right_grid_left_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_3__pin_sc_in_0_(grid_io_right_10__5__undriven_left_width_0_height_0_subtile_3__pin_sc_in_0_),
		.left_width_0_height_0_subtile_3__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_3__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_3__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_3__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_3__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_3__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_4__pin_f2a_i_0_(cby_9__2__3_right_grid_left_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_4__pin_sc_in_0_(grid_io_right_10__5__undriven_left_width_0_height_0_subtile_4__pin_sc_in_0_),
		.left_width_0_height_0_subtile_4__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_4__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_4__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_4__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_4__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_4__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_5__pin_f2a_i_0_(cby_9__2__3_right_grid_left_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_5__pin_sc_in_0_(grid_io_right_10__5__undriven_left_width_0_height_0_subtile_5__pin_sc_in_0_),
		.left_width_0_height_0_subtile_5__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_5__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_5__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_5__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_5__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_5__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_6__pin_f2a_i_0_(cby_9__2__3_right_grid_left_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_6__pin_sc_in_0_(grid_io_right_10__5__undriven_left_width_0_height_0_subtile_6__pin_sc_in_0_),
		.left_width_0_height_0_subtile_6__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_6__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_6__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_6__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_6__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_6__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_7__pin_f2a_i_0_(cby_9__2__3_right_grid_left_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_7__pin_sc_in_0_(grid_io_right_10__5__undriven_left_width_0_height_0_subtile_7__pin_sc_in_0_),
		.left_width_0_height_0_subtile_7__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_7__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_7__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_7__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_7__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_7__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_8__pin_f2a_i_0_(cby_9__2__3_right_grid_left_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_8__pin_sc_in_0_(grid_io_right_10__5__undriven_left_width_0_height_0_subtile_8__pin_sc_in_0_),
		.left_width_0_height_0_subtile_8__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_8__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_8__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_8__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_8__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_8__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_9__pin_f2a_i_0_(cby_9__2__3_right_grid_left_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_9__pin_sc_in_0_(grid_io_right_10__5__undriven_left_width_0_height_0_subtile_9__pin_sc_in_0_),
		.left_width_0_height_0_subtile_9__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_9__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_9__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_9__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_9__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_9__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_10__pin_f2a_i_0_(cby_9__2__3_right_grid_left_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_10__pin_sc_in_0_(grid_io_right_10__5__undriven_left_width_0_height_0_subtile_10__pin_sc_in_0_),
		.left_width_0_height_0_subtile_10__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_10__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_10__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_10__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_10__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_10__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_11__pin_f2a_i_0_(cby_9__2__3_right_grid_left_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_11__pin_sc_in_0_(grid_io_right_10__5__undriven_left_width_0_height_0_subtile_11__pin_sc_in_0_),
		.left_width_0_height_0_subtile_11__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_11__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_11__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_11__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_11__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_11__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_12__pin_f2a_i_0_(cby_9__2__3_right_grid_left_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_12__pin_sc_in_0_(grid_io_right_10__5__undriven_left_width_0_height_0_subtile_12__pin_sc_in_0_),
		.left_width_0_height_0_subtile_12__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_12__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_12__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_12__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_12__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_12__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_13__pin_f2a_i_0_(cby_9__2__3_right_grid_left_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_13__pin_sc_in_0_(grid_io_right_10__5__undriven_left_width_0_height_0_subtile_13__pin_sc_in_0_),
		.left_width_0_height_0_subtile_13__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_13__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_13__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_13__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_13__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_13__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_14__pin_f2a_i_0_(cby_9__2__3_right_grid_left_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_14__pin_sc_in_0_(grid_io_right_10__5__undriven_left_width_0_height_0_subtile_14__pin_sc_in_0_),
		.left_width_0_height_0_subtile_14__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_14__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_14__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_14__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_14__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_14__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_15__pin_f2a_i_0_(cby_9__2__3_right_grid_left_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_15__pin_sc_in_0_(grid_io_right_10__5__undriven_left_width_0_height_0_subtile_15__pin_sc_in_0_),
		.left_width_0_height_0_subtile_15__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_15__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_15__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_15__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_15__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_15__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_16__pin_f2a_i_0_(cby_9__2__3_right_grid_left_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_16__pin_sc_in_0_(grid_io_right_10__5__undriven_left_width_0_height_0_subtile_16__pin_sc_in_0_),
		.left_width_0_height_0_subtile_16__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_16__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_16__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_16__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_16__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_16__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_17__pin_f2a_i_0_(cby_9__2__3_right_grid_left_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_17__pin_sc_in_0_(grid_io_right_10__5__undriven_left_width_0_height_0_subtile_17__pin_sc_in_0_),
		.left_width_0_height_0_subtile_17__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_17__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_17__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_17__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_17__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_17__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_18__pin_f2a_i_0_(cby_9__2__3_right_grid_left_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_18__pin_sc_in_0_(grid_io_right_10__5__undriven_left_width_0_height_0_subtile_18__pin_sc_in_0_),
		.left_width_0_height_0_subtile_18__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_18__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_18__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_18__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_18__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_18__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_19__pin_f2a_i_0_(cby_9__2__3_right_grid_left_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_19__pin_sc_in_0_(grid_io_right_10__5__undriven_left_width_0_height_0_subtile_19__pin_sc_in_0_),
		.left_width_0_height_0_subtile_19__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_19__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_19__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_19__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_19__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_19__pin_clk_3_(clk[3]),
		.ccff_head(sb_10__1__3_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_0__pin_sc_out_0_(grid_io_right_10__5__undriven_left_width_0_height_0_subtile_0__pin_sc_out_0_),
		.left_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_1__pin_sc_out_0_(grid_io_right_10__5__undriven_left_width_0_height_0_subtile_1__pin_sc_out_0_),
		.left_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_2__pin_sc_out_0_(grid_io_right_10__5__undriven_left_width_0_height_0_subtile_2__pin_sc_out_0_),
		.left_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_3__pin_sc_out_0_(grid_io_right_10__5__undriven_left_width_0_height_0_subtile_3__pin_sc_out_0_),
		.left_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_4__pin_sc_out_0_(grid_io_right_10__5__undriven_left_width_0_height_0_subtile_4__pin_sc_out_0_),
		.left_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_5__pin_sc_out_0_(grid_io_right_10__5__undriven_left_width_0_height_0_subtile_5__pin_sc_out_0_),
		.left_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_6__pin_sc_out_0_(grid_io_right_10__5__undriven_left_width_0_height_0_subtile_6__pin_sc_out_0_),
		.left_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_7__pin_sc_out_0_(grid_io_right_10__5__undriven_left_width_0_height_0_subtile_7__pin_sc_out_0_),
		.left_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_8__pin_sc_out_0_(grid_io_right_10__5__undriven_left_width_0_height_0_subtile_8__pin_sc_out_0_),
		.left_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_9__pin_sc_out_0_(grid_io_right_10__5__undriven_left_width_0_height_0_subtile_9__pin_sc_out_0_),
		.left_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_10__pin_sc_out_0_(grid_io_right_10__5__undriven_left_width_0_height_0_subtile_10__pin_sc_out_0_),
		.left_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_11__pin_sc_out_0_(grid_io_right_10__5__undriven_left_width_0_height_0_subtile_11__pin_sc_out_0_),
		.left_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_12__pin_sc_out_0_(grid_io_right_10__5__undriven_left_width_0_height_0_subtile_12__pin_sc_out_0_),
		.left_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_13__pin_sc_out_0_(grid_io_right_10__5__undriven_left_width_0_height_0_subtile_13__pin_sc_out_0_),
		.left_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_14__pin_sc_out_0_(grid_io_right_10__5__undriven_left_width_0_height_0_subtile_14__pin_sc_out_0_),
		.left_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_15__pin_sc_out_0_(grid_io_right_10__5__undriven_left_width_0_height_0_subtile_15__pin_sc_out_0_),
		.left_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_16__pin_sc_out_0_(grid_io_right_10__5__undriven_left_width_0_height_0_subtile_16__pin_sc_out_0_),
		.left_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_17__pin_sc_out_0_(grid_io_right_10__5__undriven_left_width_0_height_0_subtile_17__pin_sc_out_0_),
		.left_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_18__pin_sc_out_0_(grid_io_right_10__5__undriven_left_width_0_height_0_subtile_18__pin_sc_out_0_),
		.left_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_19__pin_sc_out_0_(grid_io_right_10__5__undriven_left_width_0_height_0_subtile_19__pin_sc_out_0_),
		.ccff_tail(grid_io_right_4_ccff_tail));

	grid_io_right grid_io_right_10__6_ (
		.test_en(test_en),
		.scan_mode(scan_mode),
		.scan_clk(scan_clk),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.CFG_DONE(CFG_DONE),
		.gfpga_pad_QL_PREIO_A2F(gfpga_pad_QL_PREIO_A2F[360:379]),
		.gfpga_pad_QL_PREIO_F2A(gfpga_pad_QL_PREIO_F2A[360:379]),
		.gfpga_pad_QL_PREIO_F2A_DEF0(gfpga_pad_QL_PREIO_F2A_DEF0[360:379]),
		.gfpga_pad_QL_PREIO_F2A_DEF1(gfpga_pad_QL_PREIO_F2A_DEF1[360:379]),
		.gfpga_pad_QL_PREIO_F2A_CLK(gfpga_pad_QL_PREIO_F2A_CLK[360:379]),
		.left_width_0_height_0_subtile_0__pin_f2a_i_0_(cby_9__2__4_right_grid_left_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_0__pin_sc_in_0_(grid_io_right_10__6__undriven_left_width_0_height_0_subtile_0__pin_sc_in_0_),
		.left_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_1__pin_f2a_i_0_(cby_9__2__4_right_grid_left_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_1__pin_sc_in_0_(grid_io_right_10__6__undriven_left_width_0_height_0_subtile_1__pin_sc_in_0_),
		.left_width_0_height_0_subtile_1__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_1__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_1__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_1__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_1__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_1__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_2__pin_f2a_i_0_(cby_9__2__4_right_grid_left_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_2__pin_sc_in_0_(grid_io_right_10__6__undriven_left_width_0_height_0_subtile_2__pin_sc_in_0_),
		.left_width_0_height_0_subtile_2__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_2__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_2__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_2__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_2__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_2__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_3__pin_f2a_i_0_(cby_9__2__4_right_grid_left_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_3__pin_sc_in_0_(grid_io_right_10__6__undriven_left_width_0_height_0_subtile_3__pin_sc_in_0_),
		.left_width_0_height_0_subtile_3__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_3__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_3__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_3__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_3__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_3__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_4__pin_f2a_i_0_(cby_9__2__4_right_grid_left_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_4__pin_sc_in_0_(grid_io_right_10__6__undriven_left_width_0_height_0_subtile_4__pin_sc_in_0_),
		.left_width_0_height_0_subtile_4__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_4__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_4__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_4__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_4__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_4__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_5__pin_f2a_i_0_(cby_9__2__4_right_grid_left_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_5__pin_sc_in_0_(grid_io_right_10__6__undriven_left_width_0_height_0_subtile_5__pin_sc_in_0_),
		.left_width_0_height_0_subtile_5__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_5__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_5__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_5__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_5__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_5__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_6__pin_f2a_i_0_(cby_9__2__4_right_grid_left_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_6__pin_sc_in_0_(grid_io_right_10__6__undriven_left_width_0_height_0_subtile_6__pin_sc_in_0_),
		.left_width_0_height_0_subtile_6__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_6__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_6__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_6__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_6__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_6__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_7__pin_f2a_i_0_(cby_9__2__4_right_grid_left_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_7__pin_sc_in_0_(grid_io_right_10__6__undriven_left_width_0_height_0_subtile_7__pin_sc_in_0_),
		.left_width_0_height_0_subtile_7__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_7__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_7__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_7__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_7__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_7__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_8__pin_f2a_i_0_(cby_9__2__4_right_grid_left_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_8__pin_sc_in_0_(grid_io_right_10__6__undriven_left_width_0_height_0_subtile_8__pin_sc_in_0_),
		.left_width_0_height_0_subtile_8__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_8__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_8__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_8__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_8__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_8__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_9__pin_f2a_i_0_(cby_9__2__4_right_grid_left_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_9__pin_sc_in_0_(grid_io_right_10__6__undriven_left_width_0_height_0_subtile_9__pin_sc_in_0_),
		.left_width_0_height_0_subtile_9__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_9__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_9__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_9__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_9__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_9__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_10__pin_f2a_i_0_(cby_9__2__4_right_grid_left_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_10__pin_sc_in_0_(grid_io_right_10__6__undriven_left_width_0_height_0_subtile_10__pin_sc_in_0_),
		.left_width_0_height_0_subtile_10__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_10__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_10__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_10__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_10__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_10__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_11__pin_f2a_i_0_(cby_9__2__4_right_grid_left_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_11__pin_sc_in_0_(grid_io_right_10__6__undriven_left_width_0_height_0_subtile_11__pin_sc_in_0_),
		.left_width_0_height_0_subtile_11__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_11__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_11__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_11__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_11__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_11__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_12__pin_f2a_i_0_(cby_9__2__4_right_grid_left_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_12__pin_sc_in_0_(grid_io_right_10__6__undriven_left_width_0_height_0_subtile_12__pin_sc_in_0_),
		.left_width_0_height_0_subtile_12__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_12__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_12__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_12__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_12__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_12__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_13__pin_f2a_i_0_(cby_9__2__4_right_grid_left_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_13__pin_sc_in_0_(grid_io_right_10__6__undriven_left_width_0_height_0_subtile_13__pin_sc_in_0_),
		.left_width_0_height_0_subtile_13__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_13__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_13__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_13__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_13__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_13__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_14__pin_f2a_i_0_(cby_9__2__4_right_grid_left_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_14__pin_sc_in_0_(grid_io_right_10__6__undriven_left_width_0_height_0_subtile_14__pin_sc_in_0_),
		.left_width_0_height_0_subtile_14__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_14__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_14__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_14__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_14__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_14__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_15__pin_f2a_i_0_(cby_9__2__4_right_grid_left_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_15__pin_sc_in_0_(grid_io_right_10__6__undriven_left_width_0_height_0_subtile_15__pin_sc_in_0_),
		.left_width_0_height_0_subtile_15__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_15__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_15__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_15__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_15__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_15__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_16__pin_f2a_i_0_(cby_9__2__4_right_grid_left_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_16__pin_sc_in_0_(grid_io_right_10__6__undriven_left_width_0_height_0_subtile_16__pin_sc_in_0_),
		.left_width_0_height_0_subtile_16__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_16__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_16__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_16__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_16__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_16__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_17__pin_f2a_i_0_(cby_9__2__4_right_grid_left_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_17__pin_sc_in_0_(grid_io_right_10__6__undriven_left_width_0_height_0_subtile_17__pin_sc_in_0_),
		.left_width_0_height_0_subtile_17__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_17__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_17__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_17__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_17__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_17__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_18__pin_f2a_i_0_(cby_9__2__4_right_grid_left_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_18__pin_sc_in_0_(grid_io_right_10__6__undriven_left_width_0_height_0_subtile_18__pin_sc_in_0_),
		.left_width_0_height_0_subtile_18__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_18__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_18__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_18__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_18__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_18__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_19__pin_f2a_i_0_(cby_9__2__4_right_grid_left_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_19__pin_sc_in_0_(grid_io_right_10__6__undriven_left_width_0_height_0_subtile_19__pin_sc_in_0_),
		.left_width_0_height_0_subtile_19__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_19__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_19__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_19__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_19__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_19__pin_clk_3_(clk[3]),
		.ccff_head(sb_10__1__4_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_0__pin_sc_out_0_(grid_io_right_10__6__undriven_left_width_0_height_0_subtile_0__pin_sc_out_0_),
		.left_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_1__pin_sc_out_0_(grid_io_right_10__6__undriven_left_width_0_height_0_subtile_1__pin_sc_out_0_),
		.left_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_2__pin_sc_out_0_(grid_io_right_10__6__undriven_left_width_0_height_0_subtile_2__pin_sc_out_0_),
		.left_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_3__pin_sc_out_0_(grid_io_right_10__6__undriven_left_width_0_height_0_subtile_3__pin_sc_out_0_),
		.left_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_4__pin_sc_out_0_(grid_io_right_10__6__undriven_left_width_0_height_0_subtile_4__pin_sc_out_0_),
		.left_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_5__pin_sc_out_0_(grid_io_right_10__6__undriven_left_width_0_height_0_subtile_5__pin_sc_out_0_),
		.left_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_6__pin_sc_out_0_(grid_io_right_10__6__undriven_left_width_0_height_0_subtile_6__pin_sc_out_0_),
		.left_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_7__pin_sc_out_0_(grid_io_right_10__6__undriven_left_width_0_height_0_subtile_7__pin_sc_out_0_),
		.left_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_8__pin_sc_out_0_(grid_io_right_10__6__undriven_left_width_0_height_0_subtile_8__pin_sc_out_0_),
		.left_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_9__pin_sc_out_0_(grid_io_right_10__6__undriven_left_width_0_height_0_subtile_9__pin_sc_out_0_),
		.left_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_10__pin_sc_out_0_(grid_io_right_10__6__undriven_left_width_0_height_0_subtile_10__pin_sc_out_0_),
		.left_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_11__pin_sc_out_0_(grid_io_right_10__6__undriven_left_width_0_height_0_subtile_11__pin_sc_out_0_),
		.left_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_12__pin_sc_out_0_(grid_io_right_10__6__undriven_left_width_0_height_0_subtile_12__pin_sc_out_0_),
		.left_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_13__pin_sc_out_0_(grid_io_right_10__6__undriven_left_width_0_height_0_subtile_13__pin_sc_out_0_),
		.left_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_14__pin_sc_out_0_(grid_io_right_10__6__undriven_left_width_0_height_0_subtile_14__pin_sc_out_0_),
		.left_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_15__pin_sc_out_0_(grid_io_right_10__6__undriven_left_width_0_height_0_subtile_15__pin_sc_out_0_),
		.left_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_16__pin_sc_out_0_(grid_io_right_10__6__undriven_left_width_0_height_0_subtile_16__pin_sc_out_0_),
		.left_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_17__pin_sc_out_0_(grid_io_right_10__6__undriven_left_width_0_height_0_subtile_17__pin_sc_out_0_),
		.left_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_18__pin_sc_out_0_(grid_io_right_10__6__undriven_left_width_0_height_0_subtile_18__pin_sc_out_0_),
		.left_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_19__pin_sc_out_0_(grid_io_right_10__6__undriven_left_width_0_height_0_subtile_19__pin_sc_out_0_),
		.ccff_tail(grid_io_right_5_ccff_tail));

	grid_io_right grid_io_right_10__7_ (
		.test_en(test_en),
		.scan_mode(scan_mode),
		.scan_clk(scan_clk),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.CFG_DONE(CFG_DONE),
		.gfpga_pad_QL_PREIO_A2F(gfpga_pad_QL_PREIO_A2F[340:359]),
		.gfpga_pad_QL_PREIO_F2A(gfpga_pad_QL_PREIO_F2A[340:359]),
		.gfpga_pad_QL_PREIO_F2A_DEF0(gfpga_pad_QL_PREIO_F2A_DEF0[340:359]),
		.gfpga_pad_QL_PREIO_F2A_DEF1(gfpga_pad_QL_PREIO_F2A_DEF1[340:359]),
		.gfpga_pad_QL_PREIO_F2A_CLK(gfpga_pad_QL_PREIO_F2A_CLK[340:359]),
		.left_width_0_height_0_subtile_0__pin_f2a_i_0_(cby_9__2__5_right_grid_left_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_0__pin_sc_in_0_(grid_io_right_10__7__undriven_left_width_0_height_0_subtile_0__pin_sc_in_0_),
		.left_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_1__pin_f2a_i_0_(cby_9__2__5_right_grid_left_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_1__pin_sc_in_0_(grid_io_right_10__7__undriven_left_width_0_height_0_subtile_1__pin_sc_in_0_),
		.left_width_0_height_0_subtile_1__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_1__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_1__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_1__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_1__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_1__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_2__pin_f2a_i_0_(cby_9__2__5_right_grid_left_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_2__pin_sc_in_0_(grid_io_right_10__7__undriven_left_width_0_height_0_subtile_2__pin_sc_in_0_),
		.left_width_0_height_0_subtile_2__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_2__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_2__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_2__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_2__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_2__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_3__pin_f2a_i_0_(cby_9__2__5_right_grid_left_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_3__pin_sc_in_0_(grid_io_right_10__7__undriven_left_width_0_height_0_subtile_3__pin_sc_in_0_),
		.left_width_0_height_0_subtile_3__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_3__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_3__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_3__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_3__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_3__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_4__pin_f2a_i_0_(cby_9__2__5_right_grid_left_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_4__pin_sc_in_0_(grid_io_right_10__7__undriven_left_width_0_height_0_subtile_4__pin_sc_in_0_),
		.left_width_0_height_0_subtile_4__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_4__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_4__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_4__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_4__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_4__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_5__pin_f2a_i_0_(cby_9__2__5_right_grid_left_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_5__pin_sc_in_0_(grid_io_right_10__7__undriven_left_width_0_height_0_subtile_5__pin_sc_in_0_),
		.left_width_0_height_0_subtile_5__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_5__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_5__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_5__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_5__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_5__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_6__pin_f2a_i_0_(cby_9__2__5_right_grid_left_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_6__pin_sc_in_0_(grid_io_right_10__7__undriven_left_width_0_height_0_subtile_6__pin_sc_in_0_),
		.left_width_0_height_0_subtile_6__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_6__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_6__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_6__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_6__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_6__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_7__pin_f2a_i_0_(cby_9__2__5_right_grid_left_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_7__pin_sc_in_0_(grid_io_right_10__7__undriven_left_width_0_height_0_subtile_7__pin_sc_in_0_),
		.left_width_0_height_0_subtile_7__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_7__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_7__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_7__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_7__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_7__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_8__pin_f2a_i_0_(cby_9__2__5_right_grid_left_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_8__pin_sc_in_0_(grid_io_right_10__7__undriven_left_width_0_height_0_subtile_8__pin_sc_in_0_),
		.left_width_0_height_0_subtile_8__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_8__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_8__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_8__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_8__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_8__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_9__pin_f2a_i_0_(cby_9__2__5_right_grid_left_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_9__pin_sc_in_0_(grid_io_right_10__7__undriven_left_width_0_height_0_subtile_9__pin_sc_in_0_),
		.left_width_0_height_0_subtile_9__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_9__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_9__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_9__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_9__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_9__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_10__pin_f2a_i_0_(cby_9__2__5_right_grid_left_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_10__pin_sc_in_0_(grid_io_right_10__7__undriven_left_width_0_height_0_subtile_10__pin_sc_in_0_),
		.left_width_0_height_0_subtile_10__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_10__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_10__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_10__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_10__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_10__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_11__pin_f2a_i_0_(cby_9__2__5_right_grid_left_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_11__pin_sc_in_0_(grid_io_right_10__7__undriven_left_width_0_height_0_subtile_11__pin_sc_in_0_),
		.left_width_0_height_0_subtile_11__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_11__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_11__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_11__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_11__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_11__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_12__pin_f2a_i_0_(cby_9__2__5_right_grid_left_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_12__pin_sc_in_0_(grid_io_right_10__7__undriven_left_width_0_height_0_subtile_12__pin_sc_in_0_),
		.left_width_0_height_0_subtile_12__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_12__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_12__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_12__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_12__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_12__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_13__pin_f2a_i_0_(cby_9__2__5_right_grid_left_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_13__pin_sc_in_0_(grid_io_right_10__7__undriven_left_width_0_height_0_subtile_13__pin_sc_in_0_),
		.left_width_0_height_0_subtile_13__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_13__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_13__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_13__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_13__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_13__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_14__pin_f2a_i_0_(cby_9__2__5_right_grid_left_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_14__pin_sc_in_0_(grid_io_right_10__7__undriven_left_width_0_height_0_subtile_14__pin_sc_in_0_),
		.left_width_0_height_0_subtile_14__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_14__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_14__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_14__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_14__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_14__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_15__pin_f2a_i_0_(cby_9__2__5_right_grid_left_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_15__pin_sc_in_0_(grid_io_right_10__7__undriven_left_width_0_height_0_subtile_15__pin_sc_in_0_),
		.left_width_0_height_0_subtile_15__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_15__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_15__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_15__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_15__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_15__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_16__pin_f2a_i_0_(cby_9__2__5_right_grid_left_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_16__pin_sc_in_0_(grid_io_right_10__7__undriven_left_width_0_height_0_subtile_16__pin_sc_in_0_),
		.left_width_0_height_0_subtile_16__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_16__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_16__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_16__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_16__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_16__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_17__pin_f2a_i_0_(cby_9__2__5_right_grid_left_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_17__pin_sc_in_0_(grid_io_right_10__7__undriven_left_width_0_height_0_subtile_17__pin_sc_in_0_),
		.left_width_0_height_0_subtile_17__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_17__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_17__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_17__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_17__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_17__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_18__pin_f2a_i_0_(cby_9__2__5_right_grid_left_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_18__pin_sc_in_0_(grid_io_right_10__7__undriven_left_width_0_height_0_subtile_18__pin_sc_in_0_),
		.left_width_0_height_0_subtile_18__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_18__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_18__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_18__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_18__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_18__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_19__pin_f2a_i_0_(cby_9__2__5_right_grid_left_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_19__pin_sc_in_0_(grid_io_right_10__7__undriven_left_width_0_height_0_subtile_19__pin_sc_in_0_),
		.left_width_0_height_0_subtile_19__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_19__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_19__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_19__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_19__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_19__pin_clk_3_(clk[3]),
		.ccff_head(sb_10__1__5_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_0__pin_sc_out_0_(grid_io_right_10__7__undriven_left_width_0_height_0_subtile_0__pin_sc_out_0_),
		.left_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_1__pin_sc_out_0_(grid_io_right_10__7__undriven_left_width_0_height_0_subtile_1__pin_sc_out_0_),
		.left_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_2__pin_sc_out_0_(grid_io_right_10__7__undriven_left_width_0_height_0_subtile_2__pin_sc_out_0_),
		.left_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_3__pin_sc_out_0_(grid_io_right_10__7__undriven_left_width_0_height_0_subtile_3__pin_sc_out_0_),
		.left_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_4__pin_sc_out_0_(grid_io_right_10__7__undriven_left_width_0_height_0_subtile_4__pin_sc_out_0_),
		.left_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_5__pin_sc_out_0_(grid_io_right_10__7__undriven_left_width_0_height_0_subtile_5__pin_sc_out_0_),
		.left_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_6__pin_sc_out_0_(grid_io_right_10__7__undriven_left_width_0_height_0_subtile_6__pin_sc_out_0_),
		.left_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_7__pin_sc_out_0_(grid_io_right_10__7__undriven_left_width_0_height_0_subtile_7__pin_sc_out_0_),
		.left_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_8__pin_sc_out_0_(grid_io_right_10__7__undriven_left_width_0_height_0_subtile_8__pin_sc_out_0_),
		.left_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_9__pin_sc_out_0_(grid_io_right_10__7__undriven_left_width_0_height_0_subtile_9__pin_sc_out_0_),
		.left_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_10__pin_sc_out_0_(grid_io_right_10__7__undriven_left_width_0_height_0_subtile_10__pin_sc_out_0_),
		.left_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_11__pin_sc_out_0_(grid_io_right_10__7__undriven_left_width_0_height_0_subtile_11__pin_sc_out_0_),
		.left_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_12__pin_sc_out_0_(grid_io_right_10__7__undriven_left_width_0_height_0_subtile_12__pin_sc_out_0_),
		.left_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_13__pin_sc_out_0_(grid_io_right_10__7__undriven_left_width_0_height_0_subtile_13__pin_sc_out_0_),
		.left_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_14__pin_sc_out_0_(grid_io_right_10__7__undriven_left_width_0_height_0_subtile_14__pin_sc_out_0_),
		.left_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_15__pin_sc_out_0_(grid_io_right_10__7__undriven_left_width_0_height_0_subtile_15__pin_sc_out_0_),
		.left_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_16__pin_sc_out_0_(grid_io_right_10__7__undriven_left_width_0_height_0_subtile_16__pin_sc_out_0_),
		.left_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_17__pin_sc_out_0_(grid_io_right_10__7__undriven_left_width_0_height_0_subtile_17__pin_sc_out_0_),
		.left_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_18__pin_sc_out_0_(grid_io_right_10__7__undriven_left_width_0_height_0_subtile_18__pin_sc_out_0_),
		.left_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_19__pin_sc_out_0_(grid_io_right_10__7__undriven_left_width_0_height_0_subtile_19__pin_sc_out_0_),
		.ccff_tail(grid_io_right_6_ccff_tail));

	grid_io_right grid_io_right_10__8_ (
		.test_en(test_en),
		.scan_mode(scan_mode),
		.scan_clk(scan_clk),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.CFG_DONE(CFG_DONE),
		.gfpga_pad_QL_PREIO_A2F(gfpga_pad_QL_PREIO_A2F[320:339]),
		.gfpga_pad_QL_PREIO_F2A(gfpga_pad_QL_PREIO_F2A[320:339]),
		.gfpga_pad_QL_PREIO_F2A_DEF0(gfpga_pad_QL_PREIO_F2A_DEF0[320:339]),
		.gfpga_pad_QL_PREIO_F2A_DEF1(gfpga_pad_QL_PREIO_F2A_DEF1[320:339]),
		.gfpga_pad_QL_PREIO_F2A_CLK(gfpga_pad_QL_PREIO_F2A_CLK[320:339]),
		.left_width_0_height_0_subtile_0__pin_f2a_i_0_(cby_9__1__1_right_grid_left_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_0__pin_sc_in_0_(grid_io_right_10__8__undriven_left_width_0_height_0_subtile_0__pin_sc_in_0_),
		.left_width_0_height_0_subtile_0__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_0__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_0__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_0__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_0__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_1__pin_f2a_i_0_(cby_9__1__1_right_grid_left_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_1__pin_sc_in_0_(grid_io_right_10__8__undriven_left_width_0_height_0_subtile_1__pin_sc_in_0_),
		.left_width_0_height_0_subtile_1__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_1__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_1__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_1__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_1__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_1__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_2__pin_f2a_i_0_(cby_9__1__1_right_grid_left_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_2__pin_sc_in_0_(grid_io_right_10__8__undriven_left_width_0_height_0_subtile_2__pin_sc_in_0_),
		.left_width_0_height_0_subtile_2__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_2__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_2__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_2__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_2__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_2__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_3__pin_f2a_i_0_(cby_9__1__1_right_grid_left_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_3__pin_sc_in_0_(grid_io_right_10__8__undriven_left_width_0_height_0_subtile_3__pin_sc_in_0_),
		.left_width_0_height_0_subtile_3__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_3__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_3__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_3__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_3__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_3__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_4__pin_f2a_i_0_(cby_9__1__1_right_grid_left_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_4__pin_sc_in_0_(grid_io_right_10__8__undriven_left_width_0_height_0_subtile_4__pin_sc_in_0_),
		.left_width_0_height_0_subtile_4__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_4__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_4__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_4__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_4__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_4__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_5__pin_f2a_i_0_(cby_9__1__1_right_grid_left_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_5__pin_sc_in_0_(grid_io_right_10__8__undriven_left_width_0_height_0_subtile_5__pin_sc_in_0_),
		.left_width_0_height_0_subtile_5__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_5__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_5__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_5__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_5__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_5__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_6__pin_f2a_i_0_(cby_9__1__1_right_grid_left_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_6__pin_sc_in_0_(grid_io_right_10__8__undriven_left_width_0_height_0_subtile_6__pin_sc_in_0_),
		.left_width_0_height_0_subtile_6__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_6__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_6__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_6__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_6__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_6__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_7__pin_f2a_i_0_(cby_9__1__1_right_grid_left_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_7__pin_sc_in_0_(grid_io_right_10__8__undriven_left_width_0_height_0_subtile_7__pin_sc_in_0_),
		.left_width_0_height_0_subtile_7__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_7__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_7__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_7__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_7__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_7__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_8__pin_f2a_i_0_(cby_9__1__1_right_grid_left_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_8__pin_sc_in_0_(grid_io_right_10__8__undriven_left_width_0_height_0_subtile_8__pin_sc_in_0_),
		.left_width_0_height_0_subtile_8__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_8__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_8__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_8__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_8__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_8__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_9__pin_f2a_i_0_(cby_9__1__1_right_grid_left_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_9__pin_sc_in_0_(grid_io_right_10__8__undriven_left_width_0_height_0_subtile_9__pin_sc_in_0_),
		.left_width_0_height_0_subtile_9__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_9__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_9__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_9__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_9__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_9__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_10__pin_f2a_i_0_(cby_9__1__1_right_grid_left_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_10__pin_sc_in_0_(grid_io_right_10__8__undriven_left_width_0_height_0_subtile_10__pin_sc_in_0_),
		.left_width_0_height_0_subtile_10__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_10__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_10__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_10__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_10__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_10__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_11__pin_f2a_i_0_(cby_9__1__1_right_grid_left_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_11__pin_sc_in_0_(grid_io_right_10__8__undriven_left_width_0_height_0_subtile_11__pin_sc_in_0_),
		.left_width_0_height_0_subtile_11__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_11__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_11__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_11__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_11__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_11__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_12__pin_f2a_i_0_(cby_9__1__1_right_grid_left_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_12__pin_sc_in_0_(grid_io_right_10__8__undriven_left_width_0_height_0_subtile_12__pin_sc_in_0_),
		.left_width_0_height_0_subtile_12__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_12__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_12__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_12__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_12__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_12__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_13__pin_f2a_i_0_(cby_9__1__1_right_grid_left_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_13__pin_sc_in_0_(grid_io_right_10__8__undriven_left_width_0_height_0_subtile_13__pin_sc_in_0_),
		.left_width_0_height_0_subtile_13__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_13__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_13__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_13__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_13__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_13__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_14__pin_f2a_i_0_(cby_9__1__1_right_grid_left_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_14__pin_sc_in_0_(grid_io_right_10__8__undriven_left_width_0_height_0_subtile_14__pin_sc_in_0_),
		.left_width_0_height_0_subtile_14__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_14__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_14__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_14__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_14__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_14__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_15__pin_f2a_i_0_(cby_9__1__1_right_grid_left_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_15__pin_sc_in_0_(grid_io_right_10__8__undriven_left_width_0_height_0_subtile_15__pin_sc_in_0_),
		.left_width_0_height_0_subtile_15__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_15__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_15__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_15__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_15__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_15__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_16__pin_f2a_i_0_(cby_9__1__1_right_grid_left_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_16__pin_sc_in_0_(grid_io_right_10__8__undriven_left_width_0_height_0_subtile_16__pin_sc_in_0_),
		.left_width_0_height_0_subtile_16__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_16__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_16__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_16__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_16__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_16__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_17__pin_f2a_i_0_(cby_9__1__1_right_grid_left_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_17__pin_sc_in_0_(grid_io_right_10__8__undriven_left_width_0_height_0_subtile_17__pin_sc_in_0_),
		.left_width_0_height_0_subtile_17__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_17__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_17__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_17__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_17__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_17__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_18__pin_f2a_i_0_(cby_9__1__1_right_grid_left_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_18__pin_sc_in_0_(grid_io_right_10__8__undriven_left_width_0_height_0_subtile_18__pin_sc_in_0_),
		.left_width_0_height_0_subtile_18__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_18__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_18__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_18__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_18__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_18__pin_clk_3_(clk[3]),
		.left_width_0_height_0_subtile_19__pin_f2a_i_0_(cby_9__1__1_right_grid_left_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.left_width_0_height_0_subtile_19__pin_sc_in_0_(grid_io_right_10__8__undriven_left_width_0_height_0_subtile_19__pin_sc_in_0_),
		.left_width_0_height_0_subtile_19__pin_global_reset_0_(global_reset),
		.left_width_0_height_0_subtile_19__pin_scan_reset_0_(scan_reset),
		.left_width_0_height_0_subtile_19__pin_clk_0_(clk[0]),
		.left_width_0_height_0_subtile_19__pin_clk_1_(clk[1]),
		.left_width_0_height_0_subtile_19__pin_clk_2_(clk[2]),
		.left_width_0_height_0_subtile_19__pin_clk_3_(clk[3]),
		.ccff_head(sb_10__1__6_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_0__pin_sc_out_0_(grid_io_right_10__8__undriven_left_width_0_height_0_subtile_0__pin_sc_out_0_),
		.left_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_1__pin_sc_out_0_(grid_io_right_10__8__undriven_left_width_0_height_0_subtile_1__pin_sc_out_0_),
		.left_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_2__pin_sc_out_0_(grid_io_right_10__8__undriven_left_width_0_height_0_subtile_2__pin_sc_out_0_),
		.left_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_3__pin_sc_out_0_(grid_io_right_10__8__undriven_left_width_0_height_0_subtile_3__pin_sc_out_0_),
		.left_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_4__pin_sc_out_0_(grid_io_right_10__8__undriven_left_width_0_height_0_subtile_4__pin_sc_out_0_),
		.left_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_5__pin_sc_out_0_(grid_io_right_10__8__undriven_left_width_0_height_0_subtile_5__pin_sc_out_0_),
		.left_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_6__pin_sc_out_0_(grid_io_right_10__8__undriven_left_width_0_height_0_subtile_6__pin_sc_out_0_),
		.left_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_7__pin_sc_out_0_(grid_io_right_10__8__undriven_left_width_0_height_0_subtile_7__pin_sc_out_0_),
		.left_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_8__pin_sc_out_0_(grid_io_right_10__8__undriven_left_width_0_height_0_subtile_8__pin_sc_out_0_),
		.left_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_9__pin_sc_out_0_(grid_io_right_10__8__undriven_left_width_0_height_0_subtile_9__pin_sc_out_0_),
		.left_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_10__pin_sc_out_0_(grid_io_right_10__8__undriven_left_width_0_height_0_subtile_10__pin_sc_out_0_),
		.left_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_11__pin_sc_out_0_(grid_io_right_10__8__undriven_left_width_0_height_0_subtile_11__pin_sc_out_0_),
		.left_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_12__pin_sc_out_0_(grid_io_right_10__8__undriven_left_width_0_height_0_subtile_12__pin_sc_out_0_),
		.left_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_13__pin_sc_out_0_(grid_io_right_10__8__undriven_left_width_0_height_0_subtile_13__pin_sc_out_0_),
		.left_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_14__pin_sc_out_0_(grid_io_right_10__8__undriven_left_width_0_height_0_subtile_14__pin_sc_out_0_),
		.left_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_15__pin_sc_out_0_(grid_io_right_10__8__undriven_left_width_0_height_0_subtile_15__pin_sc_out_0_),
		.left_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_16__pin_sc_out_0_(grid_io_right_10__8__undriven_left_width_0_height_0_subtile_16__pin_sc_out_0_),
		.left_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_17__pin_sc_out_0_(grid_io_right_10__8__undriven_left_width_0_height_0_subtile_17__pin_sc_out_0_),
		.left_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_18__pin_sc_out_0_(grid_io_right_10__8__undriven_left_width_0_height_0_subtile_18__pin_sc_out_0_),
		.left_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.left_width_0_height_0_subtile_19__pin_sc_out_0_(grid_io_right_10__8__undriven_left_width_0_height_0_subtile_19__pin_sc_out_0_),
		.ccff_tail(ccff_tail[8]));

	sb_0__0_ sb_0__0_ (
		.chany_top_in(cby_0__1__0_chany_bottom_out[0:95]),
		.chanx_right_in(cbx_1__0__0_chanx_left_out[0:95]),
		.chany_top_out(sb_0__0__0_chany_top_out[0:95]),
		.chanx_right_out(sb_0__0__0_chanx_right_out[0:95]));

	sb_0__1_ sb_0__1_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_0__1__1_chany_bottom_out[0:95]),
		.chanx_right_in(cbx_1__0__1_chanx_left_out[0:95]),
		.chany_bottom_in(cby_0__1__0_chany_top_out[0:95]),
		.ccff_head(sb_0__1__1_ccff_tail),
		.chany_top_out(sb_0__1__0_chany_top_out[0:95]),
		.chanx_right_out(sb_0__1__0_chanx_right_out[0:95]),
		.chany_bottom_out(sb_0__1__0_chany_bottom_out[0:95]),
		.ccff_tail(sb_0__1__0_ccff_tail));

	sb_0__1_ sb_0__2_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_0__1__2_chany_bottom_out[0:95]),
		.chanx_right_in(cbx_1__0__2_chanx_left_out[0:95]),
		.chany_bottom_in(cby_0__1__1_chany_top_out[0:95]),
		.ccff_head(sb_0__1__2_ccff_tail),
		.chany_top_out(sb_0__1__1_chany_top_out[0:95]),
		.chanx_right_out(sb_0__1__1_chanx_right_out[0:95]),
		.chany_bottom_out(sb_0__1__1_chany_bottom_out[0:95]),
		.ccff_tail(sb_0__1__1_ccff_tail));

	sb_0__1_ sb_0__3_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_0__1__3_chany_bottom_out[0:95]),
		.chanx_right_in(cbx_1__0__3_chanx_left_out[0:95]),
		.chany_bottom_in(cby_0__1__2_chany_top_out[0:95]),
		.ccff_head(sb_0__1__3_ccff_tail),
		.chany_top_out(sb_0__1__2_chany_top_out[0:95]),
		.chanx_right_out(sb_0__1__2_chanx_right_out[0:95]),
		.chany_bottom_out(sb_0__1__2_chany_bottom_out[0:95]),
		.ccff_tail(sb_0__1__2_ccff_tail));

	sb_0__1_ sb_0__4_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_0__1__4_chany_bottom_out[0:95]),
		.chanx_right_in(cbx_1__0__4_chanx_left_out[0:95]),
		.chany_bottom_in(cby_0__1__3_chany_top_out[0:95]),
		.ccff_head(sb_0__1__4_ccff_tail),
		.chany_top_out(sb_0__1__3_chany_top_out[0:95]),
		.chanx_right_out(sb_0__1__3_chanx_right_out[0:95]),
		.chany_bottom_out(sb_0__1__3_chany_bottom_out[0:95]),
		.ccff_tail(sb_0__1__3_ccff_tail));

	sb_0__1_ sb_0__5_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_0__1__5_chany_bottom_out[0:95]),
		.chanx_right_in(cbx_1__0__5_chanx_left_out[0:95]),
		.chany_bottom_in(cby_0__1__4_chany_top_out[0:95]),
		.ccff_head(sb_0__1__5_ccff_tail),
		.chany_top_out(sb_0__1__4_chany_top_out[0:95]),
		.chanx_right_out(sb_0__1__4_chanx_right_out[0:95]),
		.chany_bottom_out(sb_0__1__4_chany_bottom_out[0:95]),
		.ccff_tail(sb_0__1__4_ccff_tail));

	sb_0__1_ sb_0__6_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_0__1__6_chany_bottom_out[0:95]),
		.chanx_right_in(cbx_1__0__6_chanx_left_out[0:95]),
		.chany_bottom_in(cby_0__1__5_chany_top_out[0:95]),
		.ccff_head(sb_0__1__6_ccff_tail),
		.chany_top_out(sb_0__1__5_chany_top_out[0:95]),
		.chanx_right_out(sb_0__1__5_chanx_right_out[0:95]),
		.chany_bottom_out(sb_0__1__5_chany_bottom_out[0:95]),
		.ccff_tail(sb_0__1__5_ccff_tail));

	sb_0__1_ sb_0__7_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_0__1__7_chany_bottom_out[0:95]),
		.chanx_right_in(cbx_1__0__7_chanx_left_out[0:95]),
		.chany_bottom_in(cby_0__1__6_chany_top_out[0:95]),
		.ccff_head(sb_1__8__0_ccff_tail),
		.chany_top_out(sb_0__1__6_chany_top_out[0:95]),
		.chanx_right_out(sb_0__1__6_chanx_right_out[0:95]),
		.chany_bottom_out(sb_0__1__6_chany_bottom_out[0:95]),
		.ccff_tail(sb_0__1__6_ccff_tail));

	sb_0__8_ sb_0__8_ (
		.chanx_right_in(cbx_1__0__8_chanx_left_out[0:95]),
		.chany_bottom_in(cby_0__1__7_chany_top_out[0:95]),
		.chanx_right_out(sb_0__8__0_chanx_right_out[0:95]),
		.chany_bottom_out(sb_0__8__0_chany_bottom_out[0:95]));

	sb_1__0_ sb_1__0_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_1__1__0_chany_bottom_out[0:95]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.chanx_right_in(cbx_1__0__9_chanx_left_out[0:95]),
		.chanx_left_in(cbx_1__0__0_chanx_right_out[0:95]),
		.ccff_head(sb_0__1__0_ccff_tail),
		.chany_top_out(sb_1__0__0_chany_top_out[0:95]),
		.chanx_right_out(sb_1__0__0_chanx_right_out[0:95]),
		.chanx_left_out(sb_1__0__0_chanx_left_out[0:95]),
		.ccff_tail(sb_1__0__0_ccff_tail));

	sb_1__0_ sb_9__0_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_9__1__0_chany_bottom_out[0:95]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.chanx_right_in(cbx_1__0__34_chanx_left_out[0:95]),
		.chanx_left_in(cbx_1__0__32_chanx_right_out[0:95]),
		.ccff_head(grid_io_bottom_6_ccff_tail),
		.chany_top_out(sb_1__0__1_chany_top_out[0:95]),
		.chanx_right_out(sb_1__0__1_chanx_right_out[0:95]),
		.chanx_left_out(sb_1__0__1_chanx_left_out[0:95]),
		.ccff_tail(sb_1__0__1_ccff_tail));

	sb_1__1_ sb_1__1_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_1__1__1_chany_bottom_out[0:95]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.chanx_right_in(cbx_2__1__0_chanx_left_out[0:95]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.chany_bottom_in(cby_1__1__0_chany_top_out[0:95]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_left_0_right_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.chanx_left_in(cbx_1__0__1_chanx_right_out[0:95]),
		.ccff_head(grid_clb_0_ccff_tail),
		.chany_top_out(sb_1__1__0_chany_top_out[0:95]),
		.chanx_right_out(sb_1__1__0_chanx_right_out[0:95]),
		.chany_bottom_out(sb_1__1__0_chany_bottom_out[0:95]),
		.chanx_left_out(sb_1__1__0_chanx_left_out[0:95]),
		.ccff_tail(sb_1__1__0_ccff_tail));

	sb_1__2_ sb_1__2_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_1__1__2_chany_bottom_out[0:95]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.chanx_right_in(cbx_2__2__0_chanx_left_out[0:95]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_9_),
		.chany_bottom_in(cby_1__1__1_chany_top_out[0:95]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_left_1_right_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.chanx_left_in(cbx_1__0__2_chanx_right_out[0:95]),
		.ccff_head(grid_io_left_1_ccff_tail),
		.chany_top_out(sb_1__2__0_chany_top_out[0:95]),
		.chanx_right_out(sb_1__2__0_chanx_right_out[0:95]),
		.chany_bottom_out(sb_1__2__0_chany_bottom_out[0:95]),
		.chanx_left_out(sb_1__2__0_chanx_left_out[0:95]),
		.ccff_tail(sb_1__2__0_ccff_tail));

	sb_1__2_ sb_1__3_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_1__1__3_chany_bottom_out[0:95]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.chanx_right_in(cbx_2__2__1_chanx_left_out[0:95]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_9_),
		.chany_bottom_in(cby_1__1__2_chany_top_out[0:95]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_left_2_right_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.chanx_left_in(cbx_1__0__3_chanx_right_out[0:95]),
		.ccff_head(grid_clb_2_ccff_tail),
		.chany_top_out(sb_1__2__1_chany_top_out[0:95]),
		.chanx_right_out(sb_1__2__1_chanx_right_out[0:95]),
		.chany_bottom_out(sb_1__2__1_chany_bottom_out[0:95]),
		.chanx_left_out(sb_1__2__1_chanx_left_out[0:95]),
		.ccff_tail(sb_1__2__1_ccff_tail));

	sb_1__2_ sb_1__4_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_1__1__4_chany_bottom_out[0:95]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.chanx_right_in(cbx_2__2__2_chanx_left_out[0:95]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_9_),
		.chany_bottom_in(cby_1__1__3_chany_top_out[0:95]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_left_3_right_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.chanx_left_in(cbx_1__0__4_chanx_right_out[0:95]),
		.ccff_head(grid_io_left_3_ccff_tail),
		.chany_top_out(sb_1__2__2_chany_top_out[0:95]),
		.chanx_right_out(sb_1__2__2_chanx_right_out[0:95]),
		.chany_bottom_out(sb_1__2__2_chany_bottom_out[0:95]),
		.chanx_left_out(sb_1__2__2_chanx_left_out[0:95]),
		.ccff_tail(sb_1__2__2_ccff_tail));

	sb_1__2_ sb_1__5_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_1__1__5_chany_bottom_out[0:95]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.chanx_right_in(cbx_2__2__3_chanx_left_out[0:95]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_9_),
		.chany_bottom_in(cby_1__1__4_chany_top_out[0:95]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_left_4_right_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.chanx_left_in(cbx_1__0__5_chanx_right_out[0:95]),
		.ccff_head(grid_clb_4_ccff_tail),
		.chany_top_out(sb_1__2__3_chany_top_out[0:95]),
		.chanx_right_out(sb_1__2__3_chanx_right_out[0:95]),
		.chany_bottom_out(sb_1__2__3_chany_bottom_out[0:95]),
		.chanx_left_out(sb_1__2__3_chanx_left_out[0:95]),
		.ccff_tail(sb_1__2__3_ccff_tail));

	sb_1__2_ sb_1__6_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_1__1__6_chany_bottom_out[0:95]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.chanx_right_in(cbx_2__2__4_chanx_left_out[0:95]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_9_),
		.chany_bottom_in(cby_1__1__5_chany_top_out[0:95]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_left_5_right_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.chanx_left_in(cbx_1__0__6_chanx_right_out[0:95]),
		.ccff_head(grid_io_left_5_ccff_tail),
		.chany_top_out(sb_1__2__4_chany_top_out[0:95]),
		.chanx_right_out(sb_1__2__4_chanx_right_out[0:95]),
		.chany_bottom_out(sb_1__2__4_chany_bottom_out[0:95]),
		.chanx_left_out(sb_1__2__4_chanx_left_out[0:95]),
		.ccff_tail(sb_1__2__4_ccff_tail));

	sb_1__7_ sb_1__7_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_1__1__7_chany_bottom_out[0:95]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.chanx_right_in(cbx_2__7__0_chanx_left_out[0:95]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_9_),
		.chany_bottom_in(cby_1__1__6_chany_top_out[0:95]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_left_6_right_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.chanx_left_in(cbx_1__0__7_chanx_right_out[0:95]),
		.ccff_head(grid_io_top_0_ccff_tail),
		.chany_top_out(sb_1__7__0_chany_top_out[0:95]),
		.chanx_right_out(sb_1__7__0_chanx_right_out[0:95]),
		.chany_bottom_out(sb_1__7__0_chany_bottom_out[0:95]),
		.chanx_left_out(sb_1__7__0_chanx_left_out[0:95]),
		.ccff_tail(sb_1__7__0_ccff_tail));

	sb_1__8_ sb_1__8_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chanx_right_in(cbx_1__0__10_chanx_left_out[0:95]),
		.chany_bottom_in(cby_1__1__7_chany_top_out[0:95]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_left_7_right_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.chanx_left_in(cbx_1__0__8_chanx_right_out[0:95]),
		.ccff_head(sb_2__8__0_ccff_tail),
		.chanx_right_out(sb_1__8__0_chanx_right_out[0:95]),
		.chany_bottom_out(sb_1__8__0_chany_bottom_out[0:95]),
		.chanx_left_out(sb_1__8__0_chanx_left_out[0:95]),
		.ccff_tail(sb_1__8__0_ccff_tail));

	sb_1__8_ sb_9__8_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chanx_right_in(cbx_1__0__42_chanx_left_out[0:95]),
		.chany_bottom_in(cby_9__1__1_chany_top_out[0:95]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.chanx_left_in(cbx_1__0__33_chanx_right_out[0:95]),
		.ccff_head(ccff_head[0]),
		.chanx_right_out(sb_1__8__1_chanx_right_out[0:95]),
		.chany_bottom_out(sb_1__8__1_chany_bottom_out[0:95]),
		.chanx_left_out(sb_1__8__1_chanx_left_out[0:95]),
		.ccff_tail(sb_1__8__1_ccff_tail));

	sb_2__0_ sb_2__0_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_0__1__8_chany_bottom_out[0:95]),
		.chanx_right_in(cbx_1__0__11_chanx_left_out[0:95]),
		.chanx_left_in(cbx_1__0__9_chanx_right_out[0:95]),
		.ccff_head(grid_io_left_0_ccff_tail),
		.chany_top_out(sb_2__0__0_chany_top_out[0:95]),
		.chanx_right_out(sb_2__0__0_chanx_right_out[0:95]),
		.chanx_left_out(sb_2__0__0_chanx_left_out[0:95]),
		.ccff_tail(sb_2__0__0_ccff_tail));

	sb_2__0_ sb_3__0_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_0__1__10_chany_bottom_out[0:95]),
		.chanx_right_in(cbx_1__0__13_chanx_left_out[0:95]),
		.chanx_left_in(cbx_1__0__11_chanx_right_out[0:95]),
		.ccff_head(grid_io_bottom_0_ccff_tail),
		.chany_top_out(sb_2__0__1_chany_top_out[0:95]),
		.chanx_right_out(sb_2__0__1_chanx_right_out[0:95]),
		.chanx_left_out(sb_2__0__1_chanx_left_out[0:95]),
		.ccff_tail(sb_2__0__1_ccff_tail));

	sb_2__0_ sb_4__0_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_0__1__12_chany_bottom_out[0:95]),
		.chanx_right_in(cbx_1__0__19_chanx_left_out[0:95]),
		.chanx_left_in(cbx_1__0__13_chanx_right_out[0:95]),
		.ccff_head(grid_io_bottom_1_ccff_tail),
		.chany_top_out(sb_2__0__2_chany_top_out[0:95]),
		.chanx_right_out(sb_2__0__2_chanx_right_out[0:95]),
		.chanx_left_out(sb_2__0__2_chanx_left_out[0:95]),
		.ccff_tail(sb_2__0__2_ccff_tail));

	sb_2__0_ sb_5__0_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_0__1__14_chany_bottom_out[0:95]),
		.chanx_right_in(cbx_1__0__21_chanx_left_out[0:95]),
		.chanx_left_in(cbx_1__0__19_chanx_right_out[0:95]),
		.ccff_head(grid_io_bottom_2_ccff_tail),
		.chany_top_out(sb_2__0__3_chany_top_out[0:95]),
		.chanx_right_out(sb_2__0__3_chanx_right_out[0:95]),
		.chanx_left_out(sb_2__0__3_chanx_left_out[0:95]),
		.ccff_tail(sb_2__0__3_ccff_tail));

	sb_2__0_ sb_6__0_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_0__1__16_chany_bottom_out[0:95]),
		.chanx_right_in(cbx_1__0__23_chanx_left_out[0:95]),
		.chanx_left_in(cbx_1__0__21_chanx_right_out[0:95]),
		.ccff_head(ccff_head[1]),
		.chany_top_out(sb_2__0__4_chany_top_out[0:95]),
		.chanx_right_out(sb_2__0__4_chanx_right_out[0:95]),
		.chanx_left_out(sb_2__0__4_chanx_left_out[0:95]),
		.ccff_tail(sb_2__0__4_ccff_tail));

	sb_2__0_ sb_7__0_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_0__1__18_chany_bottom_out[0:95]),
		.chanx_right_in(cbx_1__0__30_chanx_left_out[0:95]),
		.chanx_left_in(cbx_1__0__23_chanx_right_out[0:95]),
		.ccff_head(grid_io_bottom_4_ccff_tail),
		.chany_top_out(sb_2__0__5_chany_top_out[0:95]),
		.chanx_right_out(sb_2__0__5_chanx_right_out[0:95]),
		.chanx_left_out(sb_2__0__5_chanx_left_out[0:95]),
		.ccff_tail(sb_2__0__5_ccff_tail));

	sb_2__0_ sb_8__0_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_0__1__20_chany_bottom_out[0:95]),
		.chanx_right_in(cbx_1__0__32_chanx_left_out[0:95]),
		.chanx_left_in(cbx_1__0__30_chanx_right_out[0:95]),
		.ccff_head(grid_io_bottom_5_ccff_tail),
		.chany_top_out(sb_2__0__6_chany_top_out[0:95]),
		.chanx_right_out(sb_2__0__6_chanx_right_out[0:95]),
		.chanx_left_out(sb_2__0__6_chanx_left_out[0:95]),
		.ccff_tail(sb_2__0__6_ccff_tail));

	sb_2__1_ sb_2__1_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_2__2__0_chany_bottom_out[0:95]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_16_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_18_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_right_in(cbx_2__1__1_chanx_left_out[0:95]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.chany_bottom_in(cby_0__1__8_chany_top_out[0:95]),
		.chanx_left_in(cbx_2__1__0_chanx_right_out[0:95]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_bottom_0_top_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.ccff_head(grid_clb_6_ccff_tail),
		.chany_top_out(sb_2__1__0_chany_top_out[0:95]),
		.chanx_right_out(sb_2__1__0_chanx_right_out[0:95]),
		.chany_bottom_out(sb_2__1__0_chany_bottom_out[0:95]),
		.chanx_left_out(sb_2__1__0_chanx_left_out[0:95]),
		.ccff_tail(sb_2__1__0_ccff_tail));

	sb_2__1_ sb_5__1_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_2__2__12_chany_bottom_out[0:95]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_16_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_18_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_right_in(cbx_2__1__3_chanx_left_out[0:95]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.chany_bottom_in(cby_0__1__14_chany_top_out[0:95]),
		.chanx_left_in(cbx_2__1__2_chanx_right_out[0:95]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.ccff_head(grid_clb_18_ccff_tail),
		.chany_top_out(sb_2__1__1_chany_top_out[0:95]),
		.chanx_right_out(sb_2__1__1_chanx_right_out[0:95]),
		.chany_bottom_out(sb_2__1__1_chany_bottom_out[0:95]),
		.chanx_left_out(sb_2__1__1_chanx_left_out[0:95]),
		.ccff_tail(sb_2__1__1_ccff_tail));

	sb_2__1_ sb_6__1_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_2__2__18_chany_bottom_out[0:95]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_16_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_18_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_right_in(cbx_7__1__0_chanx_left_out[0:95]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.chany_bottom_in(cby_0__1__16_chany_top_out[0:95]),
		.chanx_left_in(cbx_2__1__3_chanx_right_out[0:95]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_bottom_4_top_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.ccff_head(grid_bram_0_ccff_tail),
		.chany_top_out(sb_2__1__2_chany_top_out[0:95]),
		.chanx_right_out(sb_2__1__2_chanx_right_out[0:95]),
		.chany_bottom_out(sb_2__1__2_chany_bottom_out[0:95]),
		.chanx_left_out(sb_2__1__2_chanx_left_out[0:95]),
		.ccff_tail(sb_2__1__2_ccff_tail));

	sb_2__1_ sb_8__1_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_2__2__24_chany_bottom_out[0:95]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_16_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_18_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_right_in(cbx_2__1__5_chanx_left_out[0:95]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.chany_bottom_in(cby_0__1__20_chany_top_out[0:95]),
		.chanx_left_in(cbx_2__1__4_chanx_right_out[0:95]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.ccff_head(grid_clb_30_ccff_tail),
		.chany_top_out(sb_2__1__3_chany_top_out[0:95]),
		.chanx_right_out(sb_2__1__3_chanx_right_out[0:95]),
		.chany_bottom_out(sb_2__1__3_chany_bottom_out[0:95]),
		.chanx_left_out(sb_2__1__3_chanx_left_out[0:95]),
		.ccff_tail(sb_2__1__3_ccff_tail));

	sb_2__2_ sb_2__2_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_2__2__1_chany_bottom_out[0:95]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_16_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_18_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_right_in(cbx_2__2__5_chanx_left_out[0:95]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_9_),
		.chany_bottom_in(cby_2__2__0_chany_top_out[0:95]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_left_in(cbx_2__2__0_chanx_right_out[0:95]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_7_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_9_),
		.ccff_head(grid_io_left_2_ccff_tail),
		.chany_top_out(sb_2__2__0_chany_top_out[0:95]),
		.chanx_right_out(sb_2__2__0_chanx_right_out[0:95]),
		.chany_bottom_out(sb_2__2__0_chany_bottom_out[0:95]),
		.chanx_left_out(sb_2__2__0_chanx_left_out[0:95]),
		.ccff_tail(sb_2__2__0_ccff_tail));

	sb_2__2_ sb_2__3_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_2__2__2_chany_bottom_out[0:95]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_16_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_18_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_right_in(cbx_2__2__6_chanx_left_out[0:95]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_9_),
		.chany_bottom_in(cby_2__2__1_chany_top_out[0:95]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_left_in(cbx_2__2__1_chanx_right_out[0:95]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_7_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_9_),
		.ccff_head(grid_clb_8_ccff_tail),
		.chany_top_out(sb_2__2__1_chany_top_out[0:95]),
		.chanx_right_out(sb_2__2__1_chanx_right_out[0:95]),
		.chany_bottom_out(sb_2__2__1_chany_bottom_out[0:95]),
		.chanx_left_out(sb_2__2__1_chanx_left_out[0:95]),
		.ccff_tail(sb_2__2__1_ccff_tail));

	sb_2__2_ sb_2__4_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_2__2__3_chany_bottom_out[0:95]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_16_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_18_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_right_in(cbx_2__2__7_chanx_left_out[0:95]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_9_),
		.chany_bottom_in(cby_2__2__2_chany_top_out[0:95]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_left_in(cbx_2__2__2_chanx_right_out[0:95]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_7_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_9_),
		.ccff_head(grid_io_left_4_ccff_tail),
		.chany_top_out(sb_2__2__2_chany_top_out[0:95]),
		.chanx_right_out(sb_2__2__2_chanx_right_out[0:95]),
		.chany_bottom_out(sb_2__2__2_chany_bottom_out[0:95]),
		.chanx_left_out(sb_2__2__2_chanx_left_out[0:95]),
		.ccff_tail(sb_2__2__2_ccff_tail));

	sb_2__2_ sb_2__5_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_2__2__4_chany_bottom_out[0:95]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_16_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_18_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_right_in(cbx_2__2__8_chanx_left_out[0:95]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_9_),
		.chany_bottom_in(cby_2__2__3_chany_top_out[0:95]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_left_in(cbx_2__2__3_chanx_right_out[0:95]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_7_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_9_),
		.ccff_head(grid_clb_10_ccff_tail),
		.chany_top_out(sb_2__2__3_chany_top_out[0:95]),
		.chanx_right_out(sb_2__2__3_chanx_right_out[0:95]),
		.chany_bottom_out(sb_2__2__3_chany_bottom_out[0:95]),
		.chanx_left_out(sb_2__2__3_chanx_left_out[0:95]),
		.ccff_tail(sb_2__2__3_ccff_tail));

	sb_2__2_ sb_2__6_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_2__2__5_chany_bottom_out[0:95]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_16_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_18_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_right_in(cbx_2__2__9_chanx_left_out[0:95]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_9_),
		.chany_bottom_in(cby_2__2__4_chany_top_out[0:95]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_left_in(cbx_2__2__4_chanx_right_out[0:95]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_7_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_9_),
		.ccff_head(grid_io_left_6_ccff_tail),
		.chany_top_out(sb_2__2__4_chany_top_out[0:95]),
		.chanx_right_out(sb_2__2__4_chanx_right_out[0:95]),
		.chany_bottom_out(sb_2__2__4_chany_bottom_out[0:95]),
		.chanx_left_out(sb_2__2__4_chanx_left_out[0:95]),
		.ccff_tail(sb_2__2__4_ccff_tail));

	sb_2__2_ sb_5__2_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_2__2__13_chany_bottom_out[0:95]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_16_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_18_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_right_in(cbx_2__2__15_chanx_left_out[0:95]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_9_),
		.chany_bottom_in(cby_2__2__12_chany_top_out[0:95]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_left_in(cbx_2__2__10_chanx_right_out[0:95]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_7_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_9_),
		.ccff_head(cby_4__3__0_ccff_tail),
		.chany_top_out(sb_2__2__5_chany_top_out[0:95]),
		.chanx_right_out(sb_2__2__5_chanx_right_out[0:95]),
		.chany_bottom_out(sb_2__2__5_chany_bottom_out[0:95]),
		.chanx_left_out(sb_2__2__5_chanx_left_out[0:95]),
		.ccff_tail(sb_2__2__5_ccff_tail));

	sb_2__2_ sb_5__3_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_2__2__14_chany_bottom_out[0:95]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_16_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_18_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_right_in(cbx_2__2__16_chanx_left_out[0:95]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_9_),
		.chany_bottom_in(cby_2__2__13_chany_top_out[0:95]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_left_in(cbx_2__2__11_chanx_right_out[0:95]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_7_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_9_),
		.ccff_head(grid_clb_20_ccff_tail),
		.chany_top_out(sb_2__2__6_chany_top_out[0:95]),
		.chanx_right_out(sb_2__2__6_chanx_right_out[0:95]),
		.chany_bottom_out(sb_2__2__6_chany_bottom_out[0:95]),
		.chanx_left_out(sb_2__2__6_chanx_left_out[0:95]),
		.ccff_tail(sb_2__2__6_ccff_tail));

	sb_2__2_ sb_5__4_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_2__2__15_chany_bottom_out[0:95]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_16_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_18_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_right_in(cbx_2__2__17_chanx_left_out[0:95]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_9_),
		.chany_bottom_in(cby_2__2__14_chany_top_out[0:95]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_left_in(cbx_2__2__12_chanx_right_out[0:95]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_7_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_9_),
		.ccff_head(grid_dsp_1_ccff_tail),
		.chany_top_out(sb_2__2__7_chany_top_out[0:95]),
		.chanx_right_out(sb_2__2__7_chanx_right_out[0:95]),
		.chany_bottom_out(sb_2__2__7_chany_bottom_out[0:95]),
		.chanx_left_out(sb_2__2__7_chanx_left_out[0:95]),
		.ccff_tail(sb_2__2__7_ccff_tail));

	sb_2__2_ sb_5__5_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_2__2__16_chany_bottom_out[0:95]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_16_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_18_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_right_in(cbx_2__2__18_chanx_left_out[0:95]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_9_),
		.chany_bottom_in(cby_2__2__15_chany_top_out[0:95]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_left_in(cbx_2__2__13_chanx_right_out[0:95]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_7_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_9_),
		.ccff_head(grid_clb_22_ccff_tail),
		.chany_top_out(sb_2__2__8_chany_top_out[0:95]),
		.chanx_right_out(sb_2__2__8_chanx_right_out[0:95]),
		.chany_bottom_out(sb_2__2__8_chany_bottom_out[0:95]),
		.chanx_left_out(sb_2__2__8_chanx_left_out[0:95]),
		.ccff_tail(sb_2__2__8_ccff_tail));

	sb_2__2_ sb_5__6_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_2__2__17_chany_bottom_out[0:95]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_16_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_18_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_right_in(cbx_2__2__19_chanx_left_out[0:95]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_9_),
		.chany_bottom_in(cby_2__2__16_chany_top_out[0:95]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_left_in(cbx_2__2__14_chanx_right_out[0:95]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_7_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_9_),
		.ccff_head(cby_4__4__1_ccff_tail),
		.chany_top_out(sb_2__2__9_chany_top_out[0:95]),
		.chanx_right_out(sb_2__2__9_chanx_right_out[0:95]),
		.chany_bottom_out(sb_2__2__9_chany_bottom_out[0:95]),
		.chanx_left_out(sb_2__2__9_chanx_left_out[0:95]),
		.ccff_tail(sb_2__2__9_ccff_tail));

	sb_2__2_ sb_8__2_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_2__2__25_chany_bottom_out[0:95]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_16_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_18_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_right_in(cbx_2__2__25_chanx_left_out[0:95]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_9_),
		.chany_bottom_in(cby_2__2__24_chany_top_out[0:95]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_left_in(cbx_2__2__20_chanx_right_out[0:95]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_7_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_9_),
		.ccff_head(cby_7__3__0_ccff_tail),
		.chany_top_out(sb_2__2__10_chany_top_out[0:95]),
		.chanx_right_out(sb_2__2__10_chanx_right_out[0:95]),
		.chany_bottom_out(sb_2__2__10_chany_bottom_out[0:95]),
		.chanx_left_out(sb_2__2__10_chanx_left_out[0:95]),
		.ccff_tail(sb_2__2__10_ccff_tail));

	sb_2__2_ sb_8__3_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_2__2__26_chany_bottom_out[0:95]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_16_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_18_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_right_in(cbx_2__2__26_chanx_left_out[0:95]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_9_),
		.chany_bottom_in(cby_2__2__25_chany_top_out[0:95]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_left_in(cbx_2__2__21_chanx_right_out[0:95]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_7_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_9_),
		.ccff_head(grid_clb_32_ccff_tail),
		.chany_top_out(sb_2__2__11_chany_top_out[0:95]),
		.chanx_right_out(sb_2__2__11_chanx_right_out[0:95]),
		.chany_bottom_out(sb_2__2__11_chany_bottom_out[0:95]),
		.chanx_left_out(sb_2__2__11_chanx_left_out[0:95]),
		.ccff_tail(sb_2__2__11_ccff_tail));

	sb_2__2_ sb_8__4_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_2__2__27_chany_bottom_out[0:95]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_16_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_18_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_right_in(cbx_2__2__27_chanx_left_out[0:95]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_9_),
		.chany_bottom_in(cby_2__2__26_chany_top_out[0:95]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_left_in(cbx_2__2__22_chanx_right_out[0:95]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_7_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_9_),
		.ccff_head(cby_7__5__0_ccff_tail),
		.chany_top_out(sb_2__2__12_chany_top_out[0:95]),
		.chanx_right_out(sb_2__2__12_chanx_right_out[0:95]),
		.chany_bottom_out(sb_2__2__12_chany_bottom_out[0:95]),
		.chanx_left_out(sb_2__2__12_chanx_left_out[0:95]),
		.ccff_tail(sb_2__2__12_ccff_tail));

	sb_2__2_ sb_8__5_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_2__2__28_chany_bottom_out[0:95]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_16_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_18_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_right_in(cbx_2__2__28_chanx_left_out[0:95]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_9_),
		.chany_bottom_in(cby_2__2__27_chany_top_out[0:95]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_left_in(cbx_2__2__23_chanx_right_out[0:95]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_7_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_9_),
		.ccff_head(grid_clb_34_ccff_tail),
		.chany_top_out(sb_2__2__13_chany_top_out[0:95]),
		.chanx_right_out(sb_2__2__13_chanx_right_out[0:95]),
		.chany_bottom_out(sb_2__2__13_chany_bottom_out[0:95]),
		.chanx_left_out(sb_2__2__13_chanx_left_out[0:95]),
		.ccff_tail(sb_2__2__13_ccff_tail));

	sb_2__2_ sb_8__6_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_2__2__29_chany_bottom_out[0:95]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_16_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_18_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_right_in(cbx_2__2__29_chanx_left_out[0:95]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_9_),
		.chany_bottom_in(cby_2__2__28_chany_top_out[0:95]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_left_in(cbx_2__2__24_chanx_right_out[0:95]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_7_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_9_),
		.ccff_head(cby_7__7__0_ccff_tail),
		.chany_top_out(sb_2__2__14_chany_top_out[0:95]),
		.chanx_right_out(sb_2__2__14_chanx_right_out[0:95]),
		.chany_bottom_out(sb_2__2__14_chany_bottom_out[0:95]),
		.chanx_left_out(sb_2__2__14_chanx_left_out[0:95]),
		.ccff_tail(sb_2__2__14_ccff_tail));

	sb_2__7_ sb_2__7_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_0__1__9_chany_bottom_out[0:95]),
		.chanx_right_in(cbx_2__7__1_chanx_left_out[0:95]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_9_),
		.chany_bottom_in(cby_2__2__5_chany_top_out[0:95]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_left_in(cbx_2__7__0_chanx_right_out[0:95]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_top_0_bottom_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_7_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_9_),
		.ccff_head(grid_io_top_1_ccff_tail),
		.chany_top_out(sb_2__7__0_chany_top_out[0:95]),
		.chanx_right_out(sb_2__7__0_chanx_right_out[0:95]),
		.chany_bottom_out(sb_2__7__0_chany_bottom_out[0:95]),
		.chanx_left_out(sb_2__7__0_chanx_left_out[0:95]),
		.ccff_tail(sb_2__7__0_ccff_tail));

	sb_2__7_ sb_5__7_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_0__1__15_chany_bottom_out[0:95]),
		.chanx_right_in(cbx_2__7__3_chanx_left_out[0:95]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_9_),
		.chany_bottom_in(cby_2__2__17_chany_top_out[0:95]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_left_in(cbx_2__7__2_chanx_right_out[0:95]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_7_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_9_),
		.ccff_head(grid_io_top_4_ccff_tail),
		.chany_top_out(sb_2__7__1_chany_top_out[0:95]),
		.chanx_right_out(sb_2__7__1_chanx_right_out[0:95]),
		.chany_bottom_out(sb_2__7__1_chany_bottom_out[0:95]),
		.chanx_left_out(sb_2__7__1_chanx_left_out[0:95]),
		.ccff_tail(sb_2__7__1_ccff_tail));

	sb_2__7_ sb_8__7_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_0__1__21_chany_bottom_out[0:95]),
		.chanx_right_in(cbx_2__7__5_chanx_left_out[0:95]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_9_),
		.chany_bottom_in(cby_2__2__29_chany_top_out[0:95]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_left_in(cbx_2__7__4_chanx_right_out[0:95]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_7_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_9_),
		.ccff_head(grid_io_top_7_ccff_tail),
		.chany_top_out(sb_2__7__2_chany_top_out[0:95]),
		.chanx_right_out(sb_2__7__2_chanx_right_out[0:95]),
		.chany_bottom_out(sb_2__7__2_chany_bottom_out[0:95]),
		.chanx_left_out(sb_2__7__2_chanx_left_out[0:95]),
		.ccff_tail(sb_2__7__2_ccff_tail));

	sb_2__8_ sb_2__8_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chanx_right_in(cbx_1__0__12_chanx_left_out[0:95]),
		.chany_bottom_in(cby_0__1__9_chany_top_out[0:95]),
		.chanx_left_in(cbx_1__0__10_chanx_right_out[0:95]),
		.ccff_head(sb_2__8__1_ccff_tail),
		.chanx_right_out(sb_2__8__0_chanx_right_out[0:95]),
		.chany_bottom_out(sb_2__8__0_chany_bottom_out[0:95]),
		.chanx_left_out(sb_2__8__0_chanx_left_out[0:95]),
		.ccff_tail(sb_2__8__0_ccff_tail));

	sb_2__8_ sb_3__8_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chanx_right_in(cbx_1__0__18_chanx_left_out[0:95]),
		.chany_bottom_in(cby_0__1__11_chany_top_out[0:95]),
		.chanx_left_in(cbx_1__0__12_chanx_right_out[0:95]),
		.ccff_head(sb_2__8__2_ccff_tail),
		.chanx_right_out(sb_2__8__1_chanx_right_out[0:95]),
		.chany_bottom_out(sb_2__8__1_chany_bottom_out[0:95]),
		.chanx_left_out(sb_2__8__1_chanx_left_out[0:95]),
		.ccff_tail(sb_2__8__1_ccff_tail));

	sb_2__8_ sb_4__8_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chanx_right_in(cbx_1__0__20_chanx_left_out[0:95]),
		.chany_bottom_in(cby_0__1__13_chany_top_out[0:95]),
		.chanx_left_in(cbx_1__0__18_chanx_right_out[0:95]),
		.ccff_head(sb_2__8__3_ccff_tail),
		.chanx_right_out(sb_2__8__2_chanx_right_out[0:95]),
		.chany_bottom_out(sb_2__8__2_chany_bottom_out[0:95]),
		.chanx_left_out(sb_2__8__2_chanx_left_out[0:95]),
		.ccff_tail(sb_2__8__2_ccff_tail));

	sb_2__8_ sb_5__8_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chanx_right_in(cbx_1__0__22_chanx_left_out[0:95]),
		.chany_bottom_in(cby_0__1__15_chany_top_out[0:95]),
		.chanx_left_in(cbx_1__0__20_chanx_right_out[0:95]),
		.ccff_head(sb_2__8__4_ccff_tail),
		.chanx_right_out(sb_2__8__3_chanx_right_out[0:95]),
		.chany_bottom_out(sb_2__8__3_chany_bottom_out[0:95]),
		.chanx_left_out(sb_2__8__3_chanx_left_out[0:95]),
		.ccff_tail(sb_2__8__3_ccff_tail));

	sb_2__8_ sb_6__8_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chanx_right_in(cbx_1__0__29_chanx_left_out[0:95]),
		.chany_bottom_in(cby_0__1__17_chany_top_out[0:95]),
		.chanx_left_in(cbx_1__0__22_chanx_right_out[0:95]),
		.ccff_head(sb_2__8__5_ccff_tail),
		.chanx_right_out(sb_2__8__4_chanx_right_out[0:95]),
		.chany_bottom_out(sb_2__8__4_chany_bottom_out[0:95]),
		.chanx_left_out(sb_2__8__4_chanx_left_out[0:95]),
		.ccff_tail(sb_2__8__4_ccff_tail));

	sb_2__8_ sb_7__8_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chanx_right_in(cbx_1__0__31_chanx_left_out[0:95]),
		.chany_bottom_in(cby_0__1__19_chany_top_out[0:95]),
		.chanx_left_in(cbx_1__0__29_chanx_right_out[0:95]),
		.ccff_head(sb_2__8__6_ccff_tail),
		.chanx_right_out(sb_2__8__5_chanx_right_out[0:95]),
		.chany_bottom_out(sb_2__8__5_chany_bottom_out[0:95]),
		.chanx_left_out(sb_2__8__5_chanx_left_out[0:95]),
		.ccff_tail(sb_2__8__5_ccff_tail));

	sb_2__8_ sb_8__8_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chanx_right_in(cbx_1__0__33_chanx_left_out[0:95]),
		.chany_bottom_in(cby_0__1__21_chany_top_out[0:95]),
		.chanx_left_in(cbx_1__0__31_chanx_right_out[0:95]),
		.ccff_head(sb_1__8__1_ccff_tail),
		.chanx_right_out(sb_2__8__6_chanx_right_out[0:95]),
		.chany_bottom_out(sb_2__8__6_chany_bottom_out[0:95]),
		.chanx_left_out(sb_2__8__6_chanx_left_out[0:95]),
		.ccff_tail(sb_2__8__6_ccff_tail));

	sb_3__1_ sb_3__1_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_2__2__6_chany_bottom_out[0:95]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_16_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_18_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_right_in(cbx_4__1__0_chanx_left_out[0:95]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_z_o_0_(grid_dsp_0_bottom_width_0_height_0_subtile_0__pin_z_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_z_o_1_(grid_dsp_0_bottom_width_0_height_0_subtile_0__pin_z_o_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_z_o_2_(grid_dsp_0_bottom_width_0_height_0_subtile_0__pin_z_o_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_z_o_3_(grid_dsp_0_bottom_width_0_height_0_subtile_0__pin_z_o_3_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_z_o_4_(grid_dsp_0_bottom_width_0_height_0_subtile_0__pin_z_o_4_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_z_o_5_(grid_dsp_0_bottom_width_0_height_0_subtile_0__pin_z_o_5_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_z_o_6_(grid_dsp_0_bottom_width_0_height_0_subtile_0__pin_z_o_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.chany_bottom_in(cby_0__1__10_chany_top_out[0:95]),
		.chanx_left_in(cbx_2__1__1_chanx_right_out[0:95]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_bottom_1_top_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.ccff_head(grid_dsp_0_ccff_tail),
		.chany_top_out(sb_3__1__0_chany_top_out[0:95]),
		.chanx_right_out(sb_3__1__0_chanx_right_out[0:95]),
		.chany_bottom_out(sb_3__1__0_chany_bottom_out[0:95]),
		.chanx_left_out(sb_3__1__0_chanx_left_out[0:95]),
		.ccff_tail(sb_3__1__0_ccff_tail));

	sb_3__2_ sb_3__2_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_2__2__7_chany_bottom_out[0:95]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_16_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_18_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_right_in(cbx_1__0__14_chanx_left_out[0:95]),
		.chany_bottom_in(cby_2__2__6_chany_top_out[0:95]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_left_in(cbx_2__2__5_chanx_right_out[0:95]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_7_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_9_),
		.ccff_head(ccff_head[3]),
		.chany_top_out(sb_3__2__0_chany_top_out[0:95]),
		.chanx_right_out(sb_3__2__0_chanx_right_out[0:95]),
		.chany_bottom_out(sb_3__2__0_chany_bottom_out[0:95]),
		.chanx_left_out(sb_3__2__0_chanx_left_out[0:95]),
		.ccff_tail(sb_3__2__0_ccff_tail));

	sb_3__2_ sb_3__3_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_2__2__8_chany_bottom_out[0:95]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_16_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_18_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_right_in(cbx_1__0__15_chanx_left_out[0:95]),
		.chany_bottom_in(cby_2__2__7_chany_top_out[0:95]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_left_in(cbx_2__2__6_chanx_right_out[0:95]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_7_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_9_),
		.ccff_head(cby_4__4__0_ccff_tail),
		.chany_top_out(sb_3__2__1_chany_top_out[0:95]),
		.chanx_right_out(sb_3__2__1_chanx_right_out[0:95]),
		.chany_bottom_out(sb_3__2__1_chany_bottom_out[0:95]),
		.chanx_left_out(sb_3__2__1_chanx_left_out[0:95]),
		.ccff_tail(sb_3__2__1_ccff_tail));

	sb_3__2_ sb_3__5_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_2__2__10_chany_bottom_out[0:95]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_16_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_18_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_right_in(cbx_1__0__16_chanx_left_out[0:95]),
		.chany_bottom_in(cby_2__2__9_chany_top_out[0:95]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_left_in(cbx_2__2__8_chanx_right_out[0:95]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_7_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_9_),
		.ccff_head(cby_4__3__1_ccff_tail),
		.chany_top_out(sb_3__2__2_chany_top_out[0:95]),
		.chanx_right_out(sb_3__2__2_chanx_right_out[0:95]),
		.chany_bottom_out(sb_3__2__2_chany_bottom_out[0:95]),
		.chanx_left_out(sb_3__2__2_chanx_left_out[0:95]),
		.ccff_tail(sb_3__2__2_ccff_tail));

	sb_3__2_ sb_3__6_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_2__2__11_chany_bottom_out[0:95]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_16_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_18_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_right_in(cbx_1__0__17_chanx_left_out[0:95]),
		.chany_bottom_in(cby_2__2__10_chany_top_out[0:95]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_left_in(cbx_2__2__9_chanx_right_out[0:95]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_7_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_9_),
		.ccff_head(grid_clb_5_ccff_tail),
		.chany_top_out(sb_3__2__3_chany_top_out[0:95]),
		.chanx_right_out(sb_3__2__3_chanx_right_out[0:95]),
		.chany_bottom_out(sb_3__2__3_chany_bottom_out[0:95]),
		.chanx_left_out(sb_3__2__3_chanx_left_out[0:95]),
		.ccff_tail(ccff_tail[7]));

	sb_3__2_ sb_6__2_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_2__2__19_chany_bottom_out[0:95]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_16_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_18_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_right_in(cbx_1__0__24_chanx_left_out[0:95]),
		.chany_bottom_in(cby_2__2__18_chany_top_out[0:95]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_left_in(cbx_2__2__15_chanx_right_out[0:95]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_7_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_9_),
		.ccff_head(grid_clb_13_ccff_tail),
		.chany_top_out(sb_3__2__4_chany_top_out[0:95]),
		.chanx_right_out(sb_3__2__4_chanx_right_out[0:95]),
		.chany_bottom_out(sb_3__2__4_chany_bottom_out[0:95]),
		.chanx_left_out(sb_3__2__4_chanx_left_out[0:95]),
		.ccff_tail(sb_3__2__4_ccff_tail));

	sb_3__2_ sb_6__3_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_2__2__20_chany_bottom_out[0:95]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_16_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_18_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_right_in(cbx_1__0__25_chanx_left_out[0:95]),
		.chany_bottom_in(cby_2__2__19_chany_top_out[0:95]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_left_in(cbx_2__2__16_chanx_right_out[0:95]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_7_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_9_),
		.ccff_head(cby_7__4__0_ccff_tail),
		.chany_top_out(sb_3__2__5_chany_top_out[0:95]),
		.chanx_right_out(sb_3__2__5_chanx_right_out[0:95]),
		.chany_bottom_out(sb_3__2__5_chany_bottom_out[0:95]),
		.chanx_left_out(sb_3__2__5_chanx_left_out[0:95]),
		.ccff_tail(sb_3__2__5_ccff_tail));

	sb_3__2_ sb_6__4_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_2__2__21_chany_bottom_out[0:95]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_16_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_18_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_right_in(cbx_1__0__26_chanx_left_out[0:95]),
		.chany_bottom_in(cby_2__2__20_chany_top_out[0:95]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_left_in(cbx_2__2__17_chanx_right_out[0:95]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_7_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_9_),
		.ccff_head(grid_clb_15_ccff_tail),
		.chany_top_out(sb_3__2__6_chany_top_out[0:95]),
		.chanx_right_out(sb_3__2__6_chanx_right_out[0:95]),
		.chany_bottom_out(sb_3__2__6_chany_bottom_out[0:95]),
		.chanx_left_out(sb_3__2__6_chanx_left_out[0:95]),
		.ccff_tail(sb_3__2__6_ccff_tail));

	sb_3__2_ sb_6__5_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_2__2__22_chany_bottom_out[0:95]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_16_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_18_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_right_in(cbx_1__0__27_chanx_left_out[0:95]),
		.chany_bottom_in(cby_2__2__21_chany_top_out[0:95]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_left_in(cbx_2__2__18_chanx_right_out[0:95]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_7_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_9_),
		.ccff_head(cby_7__6__0_ccff_tail),
		.chany_top_out(sb_3__2__7_chany_top_out[0:95]),
		.chanx_right_out(sb_3__2__7_chanx_right_out[0:95]),
		.chany_bottom_out(sb_3__2__7_chany_bottom_out[0:95]),
		.chanx_left_out(sb_3__2__7_chanx_left_out[0:95]),
		.ccff_tail(sb_3__2__7_ccff_tail));

	sb_3__2_ sb_6__6_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_2__2__23_chany_bottom_out[0:95]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_16_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_18_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_right_in(cbx_1__0__28_chanx_left_out[0:95]),
		.chany_bottom_in(cby_2__2__22_chany_top_out[0:95]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_left_in(cbx_2__2__19_chanx_right_out[0:95]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_7_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_9_),
		.ccff_head(grid_clb_17_ccff_tail),
		.chany_top_out(sb_3__2__8_chany_top_out[0:95]),
		.chanx_right_out(sb_3__2__8_chanx_right_out[0:95]),
		.chany_bottom_out(sb_3__2__8_chany_bottom_out[0:95]),
		.chanx_left_out(sb_3__2__8_chanx_left_out[0:95]),
		.ccff_tail(sb_3__2__8_ccff_tail));

	sb_3__4_ sb_3__4_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_2__2__9_chany_bottom_out[0:95]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_16_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_18_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_right_in(cbx_4__4__0_chanx_left_out[0:95]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_z_o_0_(grid_dsp_1_bottom_width_0_height_0_subtile_0__pin_z_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_z_o_1_(grid_dsp_1_bottom_width_0_height_0_subtile_0__pin_z_o_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_z_o_2_(grid_dsp_1_bottom_width_0_height_0_subtile_0__pin_z_o_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_z_o_3_(grid_dsp_1_bottom_width_0_height_0_subtile_0__pin_z_o_3_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_z_o_4_(grid_dsp_1_bottom_width_0_height_0_subtile_0__pin_z_o_4_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_z_o_5_(grid_dsp_1_bottom_width_0_height_0_subtile_0__pin_z_o_5_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_z_o_6_(grid_dsp_1_bottom_width_0_height_0_subtile_0__pin_z_o_6_),
		.chany_bottom_in(cby_2__2__8_chany_top_out[0:95]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_left_in(cbx_2__2__7_chanx_right_out[0:95]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_7_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_9_),
		.ccff_head(grid_clb_3_ccff_tail),
		.chany_top_out(sb_3__4__0_chany_top_out[0:95]),
		.chanx_right_out(sb_3__4__0_chanx_right_out[0:95]),
		.chany_bottom_out(sb_3__4__0_chany_bottom_out[0:95]),
		.chanx_left_out(sb_3__4__0_chanx_left_out[0:95]),
		.ccff_tail(sb_3__4__0_ccff_tail));

	sb_3__7_ sb_3__7_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_0__1__11_chany_bottom_out[0:95]),
		.chanx_right_in(cbx_4__7__0_chanx_left_out[0:95]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.chany_bottom_in(cby_2__2__11_chany_top_out[0:95]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_left_in(cbx_2__7__1_chanx_right_out[0:95]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_top_1_bottom_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_7_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_9_),
		.ccff_head(grid_io_top_2_ccff_tail),
		.chany_top_out(sb_3__7__0_chany_top_out[0:95]),
		.chanx_right_out(sb_3__7__0_chanx_right_out[0:95]),
		.chany_bottom_out(sb_3__7__0_chany_bottom_out[0:95]),
		.chanx_left_out(sb_3__7__0_chanx_left_out[0:95]),
		.ccff_tail(sb_3__7__0_ccff_tail));

	sb_3__7_ sb_6__7_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_0__1__17_chany_bottom_out[0:95]),
		.chanx_right_in(cbx_4__7__1_chanx_left_out[0:95]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.chany_bottom_in(cby_2__2__23_chany_top_out[0:95]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_left_in(cbx_2__7__3_chanx_right_out[0:95]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_top_4_bottom_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_7_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_9_),
		.ccff_head(grid_io_top_5_ccff_tail),
		.chany_top_out(sb_3__7__1_chany_top_out[0:95]),
		.chanx_right_out(sb_3__7__1_chanx_right_out[0:95]),
		.chany_bottom_out(sb_3__7__1_chany_bottom_out[0:95]),
		.chanx_left_out(sb_3__7__1_chanx_left_out[0:95]),
		.ccff_tail(sb_3__7__1_ccff_tail));

	sb_4__1_ sb_4__1_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_4__2__0_chany_bottom_out[0:95]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_z_o_7_(grid_dsp_0_right_width_0_height_0_subtile_0__pin_z_o_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_z_o_8_(grid_dsp_0_right_width_0_height_0_subtile_0__pin_z_o_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_z_o_9_(grid_dsp_0_right_width_0_height_0_subtile_0__pin_z_o_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_z_o_10_(grid_dsp_0_right_width_0_height_0_subtile_0__pin_z_o_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_z_o_11_(grid_dsp_0_right_width_0_height_0_subtile_0__pin_z_o_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_z_o_12_(grid_dsp_0_right_width_0_height_0_subtile_0__pin_z_o_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_z_o_13_(grid_dsp_0_right_width_0_height_0_subtile_0__pin_z_o_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_z_o_14_(grid_dsp_0_right_width_0_height_0_subtile_0__pin_z_o_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_z_o_15_(grid_dsp_0_right_width_0_height_0_subtile_0__pin_z_o_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_dly_b_o_0_(grid_dsp_0_right_width_0_height_0_subtile_0__pin_dly_b_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_dly_b_o_1_(grid_dsp_0_right_width_0_height_0_subtile_0__pin_dly_b_o_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_dly_b_o_2_(grid_dsp_0_right_width_0_height_0_subtile_0__pin_dly_b_o_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_dly_b_o_3_(grid_dsp_0_right_width_0_height_0_subtile_0__pin_dly_b_o_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_dly_b_o_4_(grid_dsp_0_right_width_0_height_0_subtile_0__pin_dly_b_o_4_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_dly_b_o_5_(grid_dsp_0_right_width_0_height_0_subtile_0__pin_dly_b_o_5_),
		.chanx_right_in(cbx_2__1__2_chanx_left_out[0:95]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_bottom_3_top_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.chany_bottom_in(cby_0__1__12_chany_top_out[0:95]),
		.chanx_left_in(cbx_4__1__0_chanx_right_out[0:95]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_z_o_0_(grid_dsp_0_bottom_width_0_height_0_subtile_0__pin_z_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_z_o_1_(grid_dsp_0_bottom_width_0_height_0_subtile_0__pin_z_o_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_z_o_2_(grid_dsp_0_bottom_width_0_height_0_subtile_0__pin_z_o_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_z_o_3_(grid_dsp_0_bottom_width_0_height_0_subtile_0__pin_z_o_3_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_z_o_4_(grid_dsp_0_bottom_width_0_height_0_subtile_0__pin_z_o_4_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_z_o_5_(grid_dsp_0_bottom_width_0_height_0_subtile_0__pin_z_o_5_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_z_o_6_(grid_dsp_0_bottom_width_0_height_0_subtile_0__pin_z_o_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_bottom_2_top_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.ccff_head(grid_clb_12_ccff_tail),
		.chany_top_out(sb_4__1__0_chany_top_out[0:95]),
		.chanx_right_out(sb_4__1__0_chanx_right_out[0:95]),
		.chany_bottom_out(sb_4__1__0_chany_bottom_out[0:95]),
		.chanx_left_out(sb_4__1__0_chanx_left_out[0:95]),
		.ccff_tail(sb_4__1__0_ccff_tail));

	sb_4__2_ sb_4__2_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_4__3__0_chany_bottom_out[0:95]),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_z_o_16_(grid_dsp_0_right_width_0_height_1_subtile_0__pin_z_o_16_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_z_o_17_(grid_dsp_0_right_width_0_height_1_subtile_0__pin_z_o_17_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_z_o_18_(grid_dsp_0_right_width_0_height_1_subtile_0__pin_z_o_18_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_z_o_19_(grid_dsp_0_right_width_0_height_1_subtile_0__pin_z_o_19_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_z_o_20_(grid_dsp_0_right_width_0_height_1_subtile_0__pin_z_o_20_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_z_o_21_(grid_dsp_0_right_width_0_height_1_subtile_0__pin_z_o_21_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_z_o_22_(grid_dsp_0_right_width_0_height_1_subtile_0__pin_z_o_22_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_z_o_23_(grid_dsp_0_right_width_0_height_1_subtile_0__pin_z_o_23_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_z_o_24_(grid_dsp_0_right_width_0_height_1_subtile_0__pin_z_o_24_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_z_o_25_(grid_dsp_0_right_width_0_height_1_subtile_0__pin_z_o_25_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_z_o_26_(grid_dsp_0_right_width_0_height_1_subtile_0__pin_z_o_26_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_dly_b_o_6_(grid_dsp_0_right_width_0_height_1_subtile_0__pin_dly_b_o_6_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_dly_b_o_7_(grid_dsp_0_right_width_0_height_1_subtile_0__pin_dly_b_o_7_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_dly_b_o_8_(grid_dsp_0_right_width_0_height_1_subtile_0__pin_dly_b_o_8_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_dly_b_o_9_(grid_dsp_0_right_width_0_height_1_subtile_0__pin_dly_b_o_9_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_dly_b_o_10_(grid_dsp_0_right_width_0_height_1_subtile_0__pin_dly_b_o_10_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_dly_b_o_11_(grid_dsp_0_right_width_0_height_1_subtile_0__pin_dly_b_o_11_),
		.chanx_right_in(cbx_2__2__10_chanx_left_out[0:95]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_9_),
		.chany_bottom_in(cby_4__2__0_chany_top_out[0:95]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_z_o_7_(grid_dsp_0_right_width_0_height_0_subtile_0__pin_z_o_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_z_o_8_(grid_dsp_0_right_width_0_height_0_subtile_0__pin_z_o_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_z_o_9_(grid_dsp_0_right_width_0_height_0_subtile_0__pin_z_o_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_z_o_10_(grid_dsp_0_right_width_0_height_0_subtile_0__pin_z_o_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_z_o_11_(grid_dsp_0_right_width_0_height_0_subtile_0__pin_z_o_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_z_o_12_(grid_dsp_0_right_width_0_height_0_subtile_0__pin_z_o_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_z_o_13_(grid_dsp_0_right_width_0_height_0_subtile_0__pin_z_o_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_z_o_14_(grid_dsp_0_right_width_0_height_0_subtile_0__pin_z_o_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_z_o_15_(grid_dsp_0_right_width_0_height_0_subtile_0__pin_z_o_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_dly_b_o_0_(grid_dsp_0_right_width_0_height_0_subtile_0__pin_dly_b_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_dly_b_o_1_(grid_dsp_0_right_width_0_height_0_subtile_0__pin_dly_b_o_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_dly_b_o_2_(grid_dsp_0_right_width_0_height_0_subtile_0__pin_dly_b_o_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_dly_b_o_3_(grid_dsp_0_right_width_0_height_0_subtile_0__pin_dly_b_o_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_dly_b_o_4_(grid_dsp_0_right_width_0_height_0_subtile_0__pin_dly_b_o_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_dly_b_o_5_(grid_dsp_0_right_width_0_height_0_subtile_0__pin_dly_b_o_5_),
		.chanx_left_in(cbx_1__0__14_chanx_right_out[0:95]),
		.ccff_head(grid_clb_7_ccff_tail),
		.chany_top_out(sb_4__2__0_chany_top_out[0:95]),
		.chanx_right_out(sb_4__2__0_chanx_right_out[0:95]),
		.chany_bottom_out(sb_4__2__0_chany_bottom_out[0:95]),
		.chanx_left_out(sb_4__2__0_chanx_left_out[0:95]),
		.ccff_tail(sb_4__2__0_ccff_tail));

	sb_4__2_ sb_4__5_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_4__3__1_chany_bottom_out[0:95]),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_z_o_16_(grid_dsp_1_right_width_0_height_1_subtile_0__pin_z_o_16_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_z_o_17_(grid_dsp_1_right_width_0_height_1_subtile_0__pin_z_o_17_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_z_o_18_(grid_dsp_1_right_width_0_height_1_subtile_0__pin_z_o_18_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_z_o_19_(grid_dsp_1_right_width_0_height_1_subtile_0__pin_z_o_19_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_z_o_20_(grid_dsp_1_right_width_0_height_1_subtile_0__pin_z_o_20_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_z_o_21_(grid_dsp_1_right_width_0_height_1_subtile_0__pin_z_o_21_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_z_o_22_(grid_dsp_1_right_width_0_height_1_subtile_0__pin_z_o_22_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_z_o_23_(grid_dsp_1_right_width_0_height_1_subtile_0__pin_z_o_23_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_z_o_24_(grid_dsp_1_right_width_0_height_1_subtile_0__pin_z_o_24_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_z_o_25_(grid_dsp_1_right_width_0_height_1_subtile_0__pin_z_o_25_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_z_o_26_(grid_dsp_1_right_width_0_height_1_subtile_0__pin_z_o_26_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_dly_b_o_6_(grid_dsp_1_right_width_0_height_1_subtile_0__pin_dly_b_o_6_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_dly_b_o_7_(grid_dsp_1_right_width_0_height_1_subtile_0__pin_dly_b_o_7_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_dly_b_o_8_(grid_dsp_1_right_width_0_height_1_subtile_0__pin_dly_b_o_8_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_dly_b_o_9_(grid_dsp_1_right_width_0_height_1_subtile_0__pin_dly_b_o_9_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_dly_b_o_10_(grid_dsp_1_right_width_0_height_1_subtile_0__pin_dly_b_o_10_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_dly_b_o_11_(grid_dsp_1_right_width_0_height_1_subtile_0__pin_dly_b_o_11_),
		.chanx_right_in(cbx_2__2__13_chanx_left_out[0:95]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_9_),
		.chany_bottom_in(cby_4__2__1_chany_top_out[0:95]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_z_o_7_(grid_dsp_1_right_width_0_height_0_subtile_0__pin_z_o_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_z_o_8_(grid_dsp_1_right_width_0_height_0_subtile_0__pin_z_o_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_z_o_9_(grid_dsp_1_right_width_0_height_0_subtile_0__pin_z_o_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_z_o_10_(grid_dsp_1_right_width_0_height_0_subtile_0__pin_z_o_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_z_o_11_(grid_dsp_1_right_width_0_height_0_subtile_0__pin_z_o_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_z_o_12_(grid_dsp_1_right_width_0_height_0_subtile_0__pin_z_o_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_z_o_13_(grid_dsp_1_right_width_0_height_0_subtile_0__pin_z_o_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_z_o_14_(grid_dsp_1_right_width_0_height_0_subtile_0__pin_z_o_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_z_o_15_(grid_dsp_1_right_width_0_height_0_subtile_0__pin_z_o_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_dly_b_o_0_(grid_dsp_1_right_width_0_height_0_subtile_0__pin_dly_b_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_dly_b_o_1_(grid_dsp_1_right_width_0_height_0_subtile_0__pin_dly_b_o_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_dly_b_o_2_(grid_dsp_1_right_width_0_height_0_subtile_0__pin_dly_b_o_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_dly_b_o_3_(grid_dsp_1_right_width_0_height_0_subtile_0__pin_dly_b_o_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_dly_b_o_4_(grid_dsp_1_right_width_0_height_0_subtile_0__pin_dly_b_o_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_dly_b_o_5_(grid_dsp_1_right_width_0_height_0_subtile_0__pin_dly_b_o_5_),
		.chanx_left_in(cbx_1__0__16_chanx_right_out[0:95]),
		.ccff_head(grid_clb_16_ccff_tail),
		.chany_top_out(sb_4__2__1_chany_top_out[0:95]),
		.chanx_right_out(sb_4__2__1_chanx_right_out[0:95]),
		.chany_bottom_out(sb_4__2__1_chany_bottom_out[0:95]),
		.chanx_left_out(sb_4__2__1_chanx_left_out[0:95]),
		.ccff_tail(sb_4__2__1_ccff_tail));

	sb_4__3_ sb_4__3_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_4__4__0_chany_bottom_out[0:95]),
		.top_left_grid_right_width_0_height_2_subtile_0__pin_z_o_27_(grid_dsp_0_right_width_0_height_2_subtile_0__pin_z_o_27_),
		.top_left_grid_right_width_0_height_2_subtile_0__pin_z_o_28_(grid_dsp_0_right_width_0_height_2_subtile_0__pin_z_o_28_),
		.top_left_grid_right_width_0_height_2_subtile_0__pin_z_o_29_(grid_dsp_0_right_width_0_height_2_subtile_0__pin_z_o_29_),
		.top_left_grid_right_width_0_height_2_subtile_0__pin_z_o_30_(grid_dsp_0_right_width_0_height_2_subtile_0__pin_z_o_30_),
		.top_left_grid_right_width_0_height_2_subtile_0__pin_z_o_31_(grid_dsp_0_right_width_0_height_2_subtile_0__pin_z_o_31_),
		.top_left_grid_right_width_0_height_2_subtile_0__pin_z_o_32_(grid_dsp_0_right_width_0_height_2_subtile_0__pin_z_o_32_),
		.top_left_grid_right_width_0_height_2_subtile_0__pin_z_o_33_(grid_dsp_0_right_width_0_height_2_subtile_0__pin_z_o_33_),
		.top_left_grid_right_width_0_height_2_subtile_0__pin_z_o_34_(grid_dsp_0_right_width_0_height_2_subtile_0__pin_z_o_34_),
		.top_left_grid_right_width_0_height_2_subtile_0__pin_z_o_35_(grid_dsp_0_right_width_0_height_2_subtile_0__pin_z_o_35_),
		.top_left_grid_right_width_0_height_2_subtile_0__pin_z_o_36_(grid_dsp_0_right_width_0_height_2_subtile_0__pin_z_o_36_),
		.top_left_grid_right_width_0_height_2_subtile_0__pin_z_o_37_(grid_dsp_0_right_width_0_height_2_subtile_0__pin_z_o_37_),
		.top_left_grid_right_width_0_height_2_subtile_0__pin_dly_b_o_12_(grid_dsp_0_right_width_0_height_2_subtile_0__pin_dly_b_o_12_),
		.top_left_grid_right_width_0_height_2_subtile_0__pin_dly_b_o_13_(grid_dsp_0_right_width_0_height_2_subtile_0__pin_dly_b_o_13_),
		.top_left_grid_right_width_0_height_2_subtile_0__pin_dly_b_o_14_(grid_dsp_0_right_width_0_height_2_subtile_0__pin_dly_b_o_14_),
		.top_left_grid_right_width_0_height_2_subtile_0__pin_dly_b_o_15_(grid_dsp_0_right_width_0_height_2_subtile_0__pin_dly_b_o_15_),
		.top_left_grid_right_width_0_height_2_subtile_0__pin_dly_b_o_16_(grid_dsp_0_right_width_0_height_2_subtile_0__pin_dly_b_o_16_),
		.top_left_grid_right_width_0_height_2_subtile_0__pin_dly_b_o_17_(grid_dsp_0_right_width_0_height_2_subtile_0__pin_dly_b_o_17_),
		.chanx_right_in(cbx_2__2__11_chanx_left_out[0:95]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_9_),
		.chany_bottom_in(cby_4__3__0_chany_top_out[0:95]),
		.bottom_left_grid_right_width_0_height_1_subtile_0__pin_z_o_16_(grid_dsp_0_right_width_0_height_1_subtile_0__pin_z_o_16_),
		.bottom_left_grid_right_width_0_height_1_subtile_0__pin_z_o_17_(grid_dsp_0_right_width_0_height_1_subtile_0__pin_z_o_17_),
		.bottom_left_grid_right_width_0_height_1_subtile_0__pin_z_o_18_(grid_dsp_0_right_width_0_height_1_subtile_0__pin_z_o_18_),
		.bottom_left_grid_right_width_0_height_1_subtile_0__pin_z_o_19_(grid_dsp_0_right_width_0_height_1_subtile_0__pin_z_o_19_),
		.bottom_left_grid_right_width_0_height_1_subtile_0__pin_z_o_20_(grid_dsp_0_right_width_0_height_1_subtile_0__pin_z_o_20_),
		.bottom_left_grid_right_width_0_height_1_subtile_0__pin_z_o_21_(grid_dsp_0_right_width_0_height_1_subtile_0__pin_z_o_21_),
		.bottom_left_grid_right_width_0_height_1_subtile_0__pin_z_o_22_(grid_dsp_0_right_width_0_height_1_subtile_0__pin_z_o_22_),
		.bottom_left_grid_right_width_0_height_1_subtile_0__pin_z_o_23_(grid_dsp_0_right_width_0_height_1_subtile_0__pin_z_o_23_),
		.bottom_left_grid_right_width_0_height_1_subtile_0__pin_z_o_24_(grid_dsp_0_right_width_0_height_1_subtile_0__pin_z_o_24_),
		.bottom_left_grid_right_width_0_height_1_subtile_0__pin_z_o_25_(grid_dsp_0_right_width_0_height_1_subtile_0__pin_z_o_25_),
		.bottom_left_grid_right_width_0_height_1_subtile_0__pin_z_o_26_(grid_dsp_0_right_width_0_height_1_subtile_0__pin_z_o_26_),
		.bottom_left_grid_right_width_0_height_1_subtile_0__pin_dly_b_o_6_(grid_dsp_0_right_width_0_height_1_subtile_0__pin_dly_b_o_6_),
		.bottom_left_grid_right_width_0_height_1_subtile_0__pin_dly_b_o_7_(grid_dsp_0_right_width_0_height_1_subtile_0__pin_dly_b_o_7_),
		.bottom_left_grid_right_width_0_height_1_subtile_0__pin_dly_b_o_8_(grid_dsp_0_right_width_0_height_1_subtile_0__pin_dly_b_o_8_),
		.bottom_left_grid_right_width_0_height_1_subtile_0__pin_dly_b_o_9_(grid_dsp_0_right_width_0_height_1_subtile_0__pin_dly_b_o_9_),
		.bottom_left_grid_right_width_0_height_1_subtile_0__pin_dly_b_o_10_(grid_dsp_0_right_width_0_height_1_subtile_0__pin_dly_b_o_10_),
		.bottom_left_grid_right_width_0_height_1_subtile_0__pin_dly_b_o_11_(grid_dsp_0_right_width_0_height_1_subtile_0__pin_dly_b_o_11_),
		.chanx_left_in(cbx_1__0__15_chanx_right_out[0:95]),
		.ccff_head(grid_clb_14_ccff_tail),
		.chany_top_out(sb_4__3__0_chany_top_out[0:95]),
		.chanx_right_out(sb_4__3__0_chanx_right_out[0:95]),
		.chany_bottom_out(sb_4__3__0_chany_bottom_out[0:95]),
		.chanx_left_out(sb_4__3__0_chanx_left_out[0:95]),
		.ccff_tail(sb_4__3__0_ccff_tail));

	sb_4__3_ sb_4__6_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_4__4__1_chany_bottom_out[0:95]),
		.top_left_grid_right_width_0_height_2_subtile_0__pin_z_o_27_(grid_dsp_1_right_width_0_height_2_subtile_0__pin_z_o_27_),
		.top_left_grid_right_width_0_height_2_subtile_0__pin_z_o_28_(grid_dsp_1_right_width_0_height_2_subtile_0__pin_z_o_28_),
		.top_left_grid_right_width_0_height_2_subtile_0__pin_z_o_29_(grid_dsp_1_right_width_0_height_2_subtile_0__pin_z_o_29_),
		.top_left_grid_right_width_0_height_2_subtile_0__pin_z_o_30_(grid_dsp_1_right_width_0_height_2_subtile_0__pin_z_o_30_),
		.top_left_grid_right_width_0_height_2_subtile_0__pin_z_o_31_(grid_dsp_1_right_width_0_height_2_subtile_0__pin_z_o_31_),
		.top_left_grid_right_width_0_height_2_subtile_0__pin_z_o_32_(grid_dsp_1_right_width_0_height_2_subtile_0__pin_z_o_32_),
		.top_left_grid_right_width_0_height_2_subtile_0__pin_z_o_33_(grid_dsp_1_right_width_0_height_2_subtile_0__pin_z_o_33_),
		.top_left_grid_right_width_0_height_2_subtile_0__pin_z_o_34_(grid_dsp_1_right_width_0_height_2_subtile_0__pin_z_o_34_),
		.top_left_grid_right_width_0_height_2_subtile_0__pin_z_o_35_(grid_dsp_1_right_width_0_height_2_subtile_0__pin_z_o_35_),
		.top_left_grid_right_width_0_height_2_subtile_0__pin_z_o_36_(grid_dsp_1_right_width_0_height_2_subtile_0__pin_z_o_36_),
		.top_left_grid_right_width_0_height_2_subtile_0__pin_z_o_37_(grid_dsp_1_right_width_0_height_2_subtile_0__pin_z_o_37_),
		.top_left_grid_right_width_0_height_2_subtile_0__pin_dly_b_o_12_(grid_dsp_1_right_width_0_height_2_subtile_0__pin_dly_b_o_12_),
		.top_left_grid_right_width_0_height_2_subtile_0__pin_dly_b_o_13_(grid_dsp_1_right_width_0_height_2_subtile_0__pin_dly_b_o_13_),
		.top_left_grid_right_width_0_height_2_subtile_0__pin_dly_b_o_14_(grid_dsp_1_right_width_0_height_2_subtile_0__pin_dly_b_o_14_),
		.top_left_grid_right_width_0_height_2_subtile_0__pin_dly_b_o_15_(grid_dsp_1_right_width_0_height_2_subtile_0__pin_dly_b_o_15_),
		.top_left_grid_right_width_0_height_2_subtile_0__pin_dly_b_o_16_(grid_dsp_1_right_width_0_height_2_subtile_0__pin_dly_b_o_16_),
		.top_left_grid_right_width_0_height_2_subtile_0__pin_dly_b_o_17_(grid_dsp_1_right_width_0_height_2_subtile_0__pin_dly_b_o_17_),
		.chanx_right_in(cbx_2__2__14_chanx_left_out[0:95]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_9_),
		.chany_bottom_in(cby_4__3__1_chany_top_out[0:95]),
		.bottom_left_grid_right_width_0_height_1_subtile_0__pin_z_o_16_(grid_dsp_1_right_width_0_height_1_subtile_0__pin_z_o_16_),
		.bottom_left_grid_right_width_0_height_1_subtile_0__pin_z_o_17_(grid_dsp_1_right_width_0_height_1_subtile_0__pin_z_o_17_),
		.bottom_left_grid_right_width_0_height_1_subtile_0__pin_z_o_18_(grid_dsp_1_right_width_0_height_1_subtile_0__pin_z_o_18_),
		.bottom_left_grid_right_width_0_height_1_subtile_0__pin_z_o_19_(grid_dsp_1_right_width_0_height_1_subtile_0__pin_z_o_19_),
		.bottom_left_grid_right_width_0_height_1_subtile_0__pin_z_o_20_(grid_dsp_1_right_width_0_height_1_subtile_0__pin_z_o_20_),
		.bottom_left_grid_right_width_0_height_1_subtile_0__pin_z_o_21_(grid_dsp_1_right_width_0_height_1_subtile_0__pin_z_o_21_),
		.bottom_left_grid_right_width_0_height_1_subtile_0__pin_z_o_22_(grid_dsp_1_right_width_0_height_1_subtile_0__pin_z_o_22_),
		.bottom_left_grid_right_width_0_height_1_subtile_0__pin_z_o_23_(grid_dsp_1_right_width_0_height_1_subtile_0__pin_z_o_23_),
		.bottom_left_grid_right_width_0_height_1_subtile_0__pin_z_o_24_(grid_dsp_1_right_width_0_height_1_subtile_0__pin_z_o_24_),
		.bottom_left_grid_right_width_0_height_1_subtile_0__pin_z_o_25_(grid_dsp_1_right_width_0_height_1_subtile_0__pin_z_o_25_),
		.bottom_left_grid_right_width_0_height_1_subtile_0__pin_z_o_26_(grid_dsp_1_right_width_0_height_1_subtile_0__pin_z_o_26_),
		.bottom_left_grid_right_width_0_height_1_subtile_0__pin_dly_b_o_6_(grid_dsp_1_right_width_0_height_1_subtile_0__pin_dly_b_o_6_),
		.bottom_left_grid_right_width_0_height_1_subtile_0__pin_dly_b_o_7_(grid_dsp_1_right_width_0_height_1_subtile_0__pin_dly_b_o_7_),
		.bottom_left_grid_right_width_0_height_1_subtile_0__pin_dly_b_o_8_(grid_dsp_1_right_width_0_height_1_subtile_0__pin_dly_b_o_8_),
		.bottom_left_grid_right_width_0_height_1_subtile_0__pin_dly_b_o_9_(grid_dsp_1_right_width_0_height_1_subtile_0__pin_dly_b_o_9_),
		.bottom_left_grid_right_width_0_height_1_subtile_0__pin_dly_b_o_10_(grid_dsp_1_right_width_0_height_1_subtile_0__pin_dly_b_o_10_),
		.bottom_left_grid_right_width_0_height_1_subtile_0__pin_dly_b_o_11_(grid_dsp_1_right_width_0_height_1_subtile_0__pin_dly_b_o_11_),
		.chanx_left_in(cbx_1__0__17_chanx_right_out[0:95]),
		.ccff_head(grid_clb_11_ccff_tail),
		.chany_top_out(sb_4__3__1_chany_top_out[0:95]),
		.chanx_right_out(sb_4__3__1_chanx_right_out[0:95]),
		.chany_bottom_out(sb_4__3__1_chany_bottom_out[0:95]),
		.chanx_left_out(sb_4__3__1_chanx_left_out[0:95]),
		.ccff_tail(sb_4__3__1_ccff_tail));

	sb_4__4_ sb_4__4_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_4__2__1_chany_bottom_out[0:95]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_z_o_7_(grid_dsp_1_right_width_0_height_0_subtile_0__pin_z_o_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_z_o_8_(grid_dsp_1_right_width_0_height_0_subtile_0__pin_z_o_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_z_o_9_(grid_dsp_1_right_width_0_height_0_subtile_0__pin_z_o_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_z_o_10_(grid_dsp_1_right_width_0_height_0_subtile_0__pin_z_o_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_z_o_11_(grid_dsp_1_right_width_0_height_0_subtile_0__pin_z_o_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_z_o_12_(grid_dsp_1_right_width_0_height_0_subtile_0__pin_z_o_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_z_o_13_(grid_dsp_1_right_width_0_height_0_subtile_0__pin_z_o_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_z_o_14_(grid_dsp_1_right_width_0_height_0_subtile_0__pin_z_o_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_z_o_15_(grid_dsp_1_right_width_0_height_0_subtile_0__pin_z_o_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_dly_b_o_0_(grid_dsp_1_right_width_0_height_0_subtile_0__pin_dly_b_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_dly_b_o_1_(grid_dsp_1_right_width_0_height_0_subtile_0__pin_dly_b_o_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_dly_b_o_2_(grid_dsp_1_right_width_0_height_0_subtile_0__pin_dly_b_o_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_dly_b_o_3_(grid_dsp_1_right_width_0_height_0_subtile_0__pin_dly_b_o_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_dly_b_o_4_(grid_dsp_1_right_width_0_height_0_subtile_0__pin_dly_b_o_4_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_dly_b_o_5_(grid_dsp_1_right_width_0_height_0_subtile_0__pin_dly_b_o_5_),
		.chanx_right_in(cbx_2__2__12_chanx_left_out[0:95]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_9_),
		.chany_bottom_in(cby_4__4__0_chany_top_out[0:95]),
		.bottom_left_grid_right_width_0_height_2_subtile_0__pin_z_o_27_(grid_dsp_0_right_width_0_height_2_subtile_0__pin_z_o_27_),
		.bottom_left_grid_right_width_0_height_2_subtile_0__pin_z_o_28_(grid_dsp_0_right_width_0_height_2_subtile_0__pin_z_o_28_),
		.bottom_left_grid_right_width_0_height_2_subtile_0__pin_z_o_29_(grid_dsp_0_right_width_0_height_2_subtile_0__pin_z_o_29_),
		.bottom_left_grid_right_width_0_height_2_subtile_0__pin_z_o_30_(grid_dsp_0_right_width_0_height_2_subtile_0__pin_z_o_30_),
		.bottom_left_grid_right_width_0_height_2_subtile_0__pin_z_o_31_(grid_dsp_0_right_width_0_height_2_subtile_0__pin_z_o_31_),
		.bottom_left_grid_right_width_0_height_2_subtile_0__pin_z_o_32_(grid_dsp_0_right_width_0_height_2_subtile_0__pin_z_o_32_),
		.bottom_left_grid_right_width_0_height_2_subtile_0__pin_z_o_33_(grid_dsp_0_right_width_0_height_2_subtile_0__pin_z_o_33_),
		.bottom_left_grid_right_width_0_height_2_subtile_0__pin_z_o_34_(grid_dsp_0_right_width_0_height_2_subtile_0__pin_z_o_34_),
		.bottom_left_grid_right_width_0_height_2_subtile_0__pin_z_o_35_(grid_dsp_0_right_width_0_height_2_subtile_0__pin_z_o_35_),
		.bottom_left_grid_right_width_0_height_2_subtile_0__pin_z_o_36_(grid_dsp_0_right_width_0_height_2_subtile_0__pin_z_o_36_),
		.bottom_left_grid_right_width_0_height_2_subtile_0__pin_z_o_37_(grid_dsp_0_right_width_0_height_2_subtile_0__pin_z_o_37_),
		.bottom_left_grid_right_width_0_height_2_subtile_0__pin_dly_b_o_12_(grid_dsp_0_right_width_0_height_2_subtile_0__pin_dly_b_o_12_),
		.bottom_left_grid_right_width_0_height_2_subtile_0__pin_dly_b_o_13_(grid_dsp_0_right_width_0_height_2_subtile_0__pin_dly_b_o_13_),
		.bottom_left_grid_right_width_0_height_2_subtile_0__pin_dly_b_o_14_(grid_dsp_0_right_width_0_height_2_subtile_0__pin_dly_b_o_14_),
		.bottom_left_grid_right_width_0_height_2_subtile_0__pin_dly_b_o_15_(grid_dsp_0_right_width_0_height_2_subtile_0__pin_dly_b_o_15_),
		.bottom_left_grid_right_width_0_height_2_subtile_0__pin_dly_b_o_16_(grid_dsp_0_right_width_0_height_2_subtile_0__pin_dly_b_o_16_),
		.bottom_left_grid_right_width_0_height_2_subtile_0__pin_dly_b_o_17_(grid_dsp_0_right_width_0_height_2_subtile_0__pin_dly_b_o_17_),
		.chanx_left_in(cbx_4__4__0_chanx_right_out[0:95]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_z_o_0_(grid_dsp_1_bottom_width_0_height_0_subtile_0__pin_z_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_z_o_1_(grid_dsp_1_bottom_width_0_height_0_subtile_0__pin_z_o_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_z_o_2_(grid_dsp_1_bottom_width_0_height_0_subtile_0__pin_z_o_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_z_o_3_(grid_dsp_1_bottom_width_0_height_0_subtile_0__pin_z_o_3_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_z_o_4_(grid_dsp_1_bottom_width_0_height_0_subtile_0__pin_z_o_4_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_z_o_5_(grid_dsp_1_bottom_width_0_height_0_subtile_0__pin_z_o_5_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_z_o_6_(grid_dsp_1_bottom_width_0_height_0_subtile_0__pin_z_o_6_),
		.ccff_head(grid_clb_9_ccff_tail),
		.chany_top_out(sb_4__4__0_chany_top_out[0:95]),
		.chanx_right_out(sb_4__4__0_chanx_right_out[0:95]),
		.chany_bottom_out(sb_4__4__0_chany_bottom_out[0:95]),
		.chanx_left_out(sb_4__4__0_chanx_left_out[0:95]),
		.ccff_tail(sb_4__4__0_ccff_tail));

	sb_4__7_ sb_4__7_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_0__1__13_chany_bottom_out[0:95]),
		.chanx_right_in(cbx_2__7__2_chanx_left_out[0:95]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_top_3_bottom_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_9_),
		.chany_bottom_in(cby_4__4__1_chany_top_out[0:95]),
		.bottom_left_grid_right_width_0_height_2_subtile_0__pin_z_o_27_(grid_dsp_1_right_width_0_height_2_subtile_0__pin_z_o_27_),
		.bottom_left_grid_right_width_0_height_2_subtile_0__pin_z_o_28_(grid_dsp_1_right_width_0_height_2_subtile_0__pin_z_o_28_),
		.bottom_left_grid_right_width_0_height_2_subtile_0__pin_z_o_29_(grid_dsp_1_right_width_0_height_2_subtile_0__pin_z_o_29_),
		.bottom_left_grid_right_width_0_height_2_subtile_0__pin_z_o_30_(grid_dsp_1_right_width_0_height_2_subtile_0__pin_z_o_30_),
		.bottom_left_grid_right_width_0_height_2_subtile_0__pin_z_o_31_(grid_dsp_1_right_width_0_height_2_subtile_0__pin_z_o_31_),
		.bottom_left_grid_right_width_0_height_2_subtile_0__pin_z_o_32_(grid_dsp_1_right_width_0_height_2_subtile_0__pin_z_o_32_),
		.bottom_left_grid_right_width_0_height_2_subtile_0__pin_z_o_33_(grid_dsp_1_right_width_0_height_2_subtile_0__pin_z_o_33_),
		.bottom_left_grid_right_width_0_height_2_subtile_0__pin_z_o_34_(grid_dsp_1_right_width_0_height_2_subtile_0__pin_z_o_34_),
		.bottom_left_grid_right_width_0_height_2_subtile_0__pin_z_o_35_(grid_dsp_1_right_width_0_height_2_subtile_0__pin_z_o_35_),
		.bottom_left_grid_right_width_0_height_2_subtile_0__pin_z_o_36_(grid_dsp_1_right_width_0_height_2_subtile_0__pin_z_o_36_),
		.bottom_left_grid_right_width_0_height_2_subtile_0__pin_z_o_37_(grid_dsp_1_right_width_0_height_2_subtile_0__pin_z_o_37_),
		.bottom_left_grid_right_width_0_height_2_subtile_0__pin_dly_b_o_12_(grid_dsp_1_right_width_0_height_2_subtile_0__pin_dly_b_o_12_),
		.bottom_left_grid_right_width_0_height_2_subtile_0__pin_dly_b_o_13_(grid_dsp_1_right_width_0_height_2_subtile_0__pin_dly_b_o_13_),
		.bottom_left_grid_right_width_0_height_2_subtile_0__pin_dly_b_o_14_(grid_dsp_1_right_width_0_height_2_subtile_0__pin_dly_b_o_14_),
		.bottom_left_grid_right_width_0_height_2_subtile_0__pin_dly_b_o_15_(grid_dsp_1_right_width_0_height_2_subtile_0__pin_dly_b_o_15_),
		.bottom_left_grid_right_width_0_height_2_subtile_0__pin_dly_b_o_16_(grid_dsp_1_right_width_0_height_2_subtile_0__pin_dly_b_o_16_),
		.bottom_left_grid_right_width_0_height_2_subtile_0__pin_dly_b_o_17_(grid_dsp_1_right_width_0_height_2_subtile_0__pin_dly_b_o_17_),
		.chanx_left_in(cbx_4__7__0_chanx_right_out[0:95]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_top_2_bottom_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.ccff_head(grid_io_top_3_ccff_tail),
		.chany_top_out(sb_4__7__0_chany_top_out[0:95]),
		.chanx_right_out(sb_4__7__0_chanx_right_out[0:95]),
		.chany_bottom_out(sb_4__7__0_chany_bottom_out[0:95]),
		.chanx_left_out(sb_4__7__0_chanx_left_out[0:95]),
		.ccff_tail(sb_4__7__0_ccff_tail));

	sb_7__1_ sb_7__1_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_7__2__0_chany_bottom_out[0:95]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_A1_o_0_(grid_bram_0_right_width_0_height_0_subtile_0__pin_RDATA_A1_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_A1_o_1_(grid_bram_0_right_width_0_height_0_subtile_0__pin_RDATA_A1_o_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_A1_o_2_(grid_bram_0_right_width_0_height_0_subtile_0__pin_RDATA_A1_o_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_A1_o_3_(grid_bram_0_right_width_0_height_0_subtile_0__pin_RDATA_A1_o_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_A1_o_4_(grid_bram_0_right_width_0_height_0_subtile_0__pin_RDATA_A1_o_4_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_A1_o_5_(grid_bram_0_right_width_0_height_0_subtile_0__pin_RDATA_A1_o_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_B1_o_0_(grid_bram_0_right_width_0_height_0_subtile_0__pin_RDATA_B1_o_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_B1_o_1_(grid_bram_0_right_width_0_height_0_subtile_0__pin_RDATA_B1_o_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_B1_o_2_(grid_bram_0_right_width_0_height_0_subtile_0__pin_RDATA_B1_o_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_B1_o_3_(grid_bram_0_right_width_0_height_0_subtile_0__pin_RDATA_B1_o_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_B1_o_4_(grid_bram_0_right_width_0_height_0_subtile_0__pin_RDATA_B1_o_4_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_B1_o_5_(grid_bram_0_right_width_0_height_0_subtile_0__pin_RDATA_B1_o_5_),
		.chanx_right_in(cbx_2__1__4_chanx_left_out[0:95]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_bottom_6_top_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.chany_bottom_in(cby_0__1__18_chany_top_out[0:95]),
		.chanx_left_in(cbx_7__1__0_chanx_right_out[0:95]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_bottom_5_top_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.ccff_head(grid_clb_24_ccff_tail),
		.chany_top_out(sb_7__1__0_chany_top_out[0:95]),
		.chanx_right_out(sb_7__1__0_chanx_right_out[0:95]),
		.chany_bottom_out(sb_7__1__0_chany_bottom_out[0:95]),
		.chanx_left_out(sb_7__1__0_chanx_left_out[0:95]),
		.ccff_tail(sb_7__1__0_ccff_tail));

	sb_7__2_ sb_7__2_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_7__3__0_chany_bottom_out[0:95]),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_A1_o_6_(grid_bram_0_right_width_0_height_1_subtile_0__pin_RDATA_A1_o_6_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_A1_o_7_(grid_bram_0_right_width_0_height_1_subtile_0__pin_RDATA_A1_o_7_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_A1_o_8_(grid_bram_0_right_width_0_height_1_subtile_0__pin_RDATA_A1_o_8_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_A1_o_9_(grid_bram_0_right_width_0_height_1_subtile_0__pin_RDATA_A1_o_9_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_A1_o_10_(grid_bram_0_right_width_0_height_1_subtile_0__pin_RDATA_A1_o_10_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_A1_o_11_(grid_bram_0_right_width_0_height_1_subtile_0__pin_RDATA_A1_o_11_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_B1_o_6_(grid_bram_0_right_width_0_height_1_subtile_0__pin_RDATA_B1_o_6_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_B1_o_7_(grid_bram_0_right_width_0_height_1_subtile_0__pin_RDATA_B1_o_7_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_B1_o_8_(grid_bram_0_right_width_0_height_1_subtile_0__pin_RDATA_B1_o_8_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_B1_o_9_(grid_bram_0_right_width_0_height_1_subtile_0__pin_RDATA_B1_o_9_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_B1_o_10_(grid_bram_0_right_width_0_height_1_subtile_0__pin_RDATA_B1_o_10_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_B1_o_11_(grid_bram_0_right_width_0_height_1_subtile_0__pin_RDATA_B1_o_11_),
		.chanx_right_in(cbx_2__2__20_chanx_left_out[0:95]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_9_),
		.chany_bottom_in(cby_7__2__0_chany_top_out[0:95]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_A1_o_0_(grid_bram_0_right_width_0_height_0_subtile_0__pin_RDATA_A1_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_A1_o_1_(grid_bram_0_right_width_0_height_0_subtile_0__pin_RDATA_A1_o_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_A1_o_2_(grid_bram_0_right_width_0_height_0_subtile_0__pin_RDATA_A1_o_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_A1_o_3_(grid_bram_0_right_width_0_height_0_subtile_0__pin_RDATA_A1_o_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_A1_o_4_(grid_bram_0_right_width_0_height_0_subtile_0__pin_RDATA_A1_o_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_A1_o_5_(grid_bram_0_right_width_0_height_0_subtile_0__pin_RDATA_A1_o_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_B1_o_0_(grid_bram_0_right_width_0_height_0_subtile_0__pin_RDATA_B1_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_B1_o_1_(grid_bram_0_right_width_0_height_0_subtile_0__pin_RDATA_B1_o_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_B1_o_2_(grid_bram_0_right_width_0_height_0_subtile_0__pin_RDATA_B1_o_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_B1_o_3_(grid_bram_0_right_width_0_height_0_subtile_0__pin_RDATA_B1_o_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_B1_o_4_(grid_bram_0_right_width_0_height_0_subtile_0__pin_RDATA_B1_o_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_B1_o_5_(grid_bram_0_right_width_0_height_0_subtile_0__pin_RDATA_B1_o_5_),
		.chanx_left_in(cbx_1__0__24_chanx_right_out[0:95]),
		.ccff_head(grid_clb_19_ccff_tail),
		.chany_top_out(sb_7__2__0_chany_top_out[0:95]),
		.chanx_right_out(sb_7__2__0_chanx_right_out[0:95]),
		.chany_bottom_out(sb_7__2__0_chany_bottom_out[0:95]),
		.chanx_left_out(sb_7__2__0_chanx_left_out[0:95]),
		.ccff_tail(sb_7__2__0_ccff_tail));

	sb_7__2_ sb_7__3_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_7__4__0_chany_bottom_out[0:95]),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_A1_o_6_(grid_bram_0_right_width_0_height_2_subtile_0__pin_RDATA_A1_o_12_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_A1_o_7_(grid_bram_0_right_width_0_height_2_subtile_0__pin_RDATA_A1_o_13_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_A1_o_8_(grid_bram_0_right_width_0_height_2_subtile_0__pin_RDATA_A1_o_14_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_A1_o_9_(grid_bram_0_right_width_0_height_2_subtile_0__pin_RDATA_A1_o_15_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_A1_o_10_(grid_bram_0_right_width_0_height_2_subtile_0__pin_RDATA_A1_o_16_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_A1_o_11_(grid_bram_0_right_width_0_height_2_subtile_0__pin_RDATA_A1_o_17_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_B1_o_6_(grid_bram_0_right_width_0_height_2_subtile_0__pin_RDATA_B1_o_12_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_B1_o_7_(grid_bram_0_right_width_0_height_2_subtile_0__pin_RDATA_B1_o_13_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_B1_o_8_(grid_bram_0_right_width_0_height_2_subtile_0__pin_RDATA_B1_o_14_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_B1_o_9_(grid_bram_0_right_width_0_height_2_subtile_0__pin_RDATA_B1_o_15_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_B1_o_10_(grid_bram_0_right_width_0_height_2_subtile_0__pin_RDATA_B1_o_16_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_B1_o_11_(grid_bram_0_right_width_0_height_2_subtile_0__pin_RDATA_B1_o_17_),
		.chanx_right_in(cbx_2__2__21_chanx_left_out[0:95]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_9_),
		.chany_bottom_in(cby_7__3__0_chany_top_out[0:95]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_A1_o_0_(grid_bram_0_right_width_0_height_1_subtile_0__pin_RDATA_A1_o_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_A1_o_1_(grid_bram_0_right_width_0_height_1_subtile_0__pin_RDATA_A1_o_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_A1_o_2_(grid_bram_0_right_width_0_height_1_subtile_0__pin_RDATA_A1_o_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_A1_o_3_(grid_bram_0_right_width_0_height_1_subtile_0__pin_RDATA_A1_o_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_A1_o_4_(grid_bram_0_right_width_0_height_1_subtile_0__pin_RDATA_A1_o_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_A1_o_5_(grid_bram_0_right_width_0_height_1_subtile_0__pin_RDATA_A1_o_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_B1_o_0_(grid_bram_0_right_width_0_height_1_subtile_0__pin_RDATA_B1_o_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_B1_o_1_(grid_bram_0_right_width_0_height_1_subtile_0__pin_RDATA_B1_o_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_B1_o_2_(grid_bram_0_right_width_0_height_1_subtile_0__pin_RDATA_B1_o_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_B1_o_3_(grid_bram_0_right_width_0_height_1_subtile_0__pin_RDATA_B1_o_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_B1_o_4_(grid_bram_0_right_width_0_height_1_subtile_0__pin_RDATA_B1_o_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_B1_o_5_(grid_bram_0_right_width_0_height_1_subtile_0__pin_RDATA_B1_o_11_),
		.chanx_left_in(cbx_1__0__25_chanx_right_out[0:95]),
		.ccff_head(grid_clb_26_ccff_tail),
		.chany_top_out(sb_7__2__1_chany_top_out[0:95]),
		.chanx_right_out(sb_7__2__1_chanx_right_out[0:95]),
		.chany_bottom_out(sb_7__2__1_chany_bottom_out[0:95]),
		.chanx_left_out(sb_7__2__1_chanx_left_out[0:95]),
		.ccff_tail(sb_7__2__1_ccff_tail));

	sb_7__2_ sb_7__4_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_7__5__0_chany_bottom_out[0:95]),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_A1_o_6_(grid_bram_0_right_width_0_height_3_subtile_0__pin_RDATA_A2_o_0_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_A1_o_7_(grid_bram_0_right_width_0_height_3_subtile_0__pin_RDATA_A2_o_1_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_A1_o_8_(grid_bram_0_right_width_0_height_3_subtile_0__pin_RDATA_A2_o_2_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_A1_o_9_(grid_bram_0_right_width_0_height_3_subtile_0__pin_RDATA_A2_o_3_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_A1_o_10_(grid_bram_0_right_width_0_height_3_subtile_0__pin_RDATA_A2_o_4_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_A1_o_11_(grid_bram_0_right_width_0_height_3_subtile_0__pin_RDATA_A2_o_5_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_B1_o_6_(grid_bram_0_right_width_0_height_3_subtile_0__pin_RDATA_B2_o_0_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_B1_o_7_(grid_bram_0_right_width_0_height_3_subtile_0__pin_RDATA_B2_o_1_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_B1_o_8_(grid_bram_0_right_width_0_height_3_subtile_0__pin_RDATA_B2_o_2_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_B1_o_9_(grid_bram_0_right_width_0_height_3_subtile_0__pin_RDATA_B2_o_3_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_B1_o_10_(grid_bram_0_right_width_0_height_3_subtile_0__pin_RDATA_B2_o_4_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_B1_o_11_(grid_bram_0_right_width_0_height_3_subtile_0__pin_RDATA_B2_o_5_),
		.chanx_right_in(cbx_2__2__22_chanx_left_out[0:95]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_9_),
		.chany_bottom_in(cby_7__4__0_chany_top_out[0:95]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_A1_o_0_(grid_bram_0_right_width_0_height_2_subtile_0__pin_RDATA_A1_o_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_A1_o_1_(grid_bram_0_right_width_0_height_2_subtile_0__pin_RDATA_A1_o_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_A1_o_2_(grid_bram_0_right_width_0_height_2_subtile_0__pin_RDATA_A1_o_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_A1_o_3_(grid_bram_0_right_width_0_height_2_subtile_0__pin_RDATA_A1_o_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_A1_o_4_(grid_bram_0_right_width_0_height_2_subtile_0__pin_RDATA_A1_o_16_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_A1_o_5_(grid_bram_0_right_width_0_height_2_subtile_0__pin_RDATA_A1_o_17_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_B1_o_0_(grid_bram_0_right_width_0_height_2_subtile_0__pin_RDATA_B1_o_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_B1_o_1_(grid_bram_0_right_width_0_height_2_subtile_0__pin_RDATA_B1_o_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_B1_o_2_(grid_bram_0_right_width_0_height_2_subtile_0__pin_RDATA_B1_o_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_B1_o_3_(grid_bram_0_right_width_0_height_2_subtile_0__pin_RDATA_B1_o_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_B1_o_4_(grid_bram_0_right_width_0_height_2_subtile_0__pin_RDATA_B1_o_16_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_B1_o_5_(grid_bram_0_right_width_0_height_2_subtile_0__pin_RDATA_B1_o_17_),
		.chanx_left_in(cbx_1__0__26_chanx_right_out[0:95]),
		.ccff_head(grid_clb_21_ccff_tail),
		.chany_top_out(sb_7__2__2_chany_top_out[0:95]),
		.chanx_right_out(sb_7__2__2_chanx_right_out[0:95]),
		.chany_bottom_out(sb_7__2__2_chany_bottom_out[0:95]),
		.chanx_left_out(sb_7__2__2_chanx_left_out[0:95]),
		.ccff_tail(sb_7__2__2_ccff_tail));

	sb_7__2_ sb_7__5_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_7__6__0_chany_bottom_out[0:95]),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_A1_o_6_(grid_bram_0_right_width_0_height_4_subtile_0__pin_RDATA_A2_o_6_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_A1_o_7_(grid_bram_0_right_width_0_height_4_subtile_0__pin_RDATA_A2_o_7_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_A1_o_8_(grid_bram_0_right_width_0_height_4_subtile_0__pin_RDATA_A2_o_8_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_A1_o_9_(grid_bram_0_right_width_0_height_4_subtile_0__pin_RDATA_A2_o_9_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_A1_o_10_(grid_bram_0_right_width_0_height_4_subtile_0__pin_RDATA_A2_o_10_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_A1_o_11_(grid_bram_0_right_width_0_height_4_subtile_0__pin_RDATA_A2_o_11_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_B1_o_6_(grid_bram_0_right_width_0_height_4_subtile_0__pin_RDATA_B2_o_6_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_B1_o_7_(grid_bram_0_right_width_0_height_4_subtile_0__pin_RDATA_B2_o_7_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_B1_o_8_(grid_bram_0_right_width_0_height_4_subtile_0__pin_RDATA_B2_o_8_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_B1_o_9_(grid_bram_0_right_width_0_height_4_subtile_0__pin_RDATA_B2_o_9_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_B1_o_10_(grid_bram_0_right_width_0_height_4_subtile_0__pin_RDATA_B2_o_10_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_B1_o_11_(grid_bram_0_right_width_0_height_4_subtile_0__pin_RDATA_B2_o_11_),
		.chanx_right_in(cbx_2__2__23_chanx_left_out[0:95]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_9_),
		.chany_bottom_in(cby_7__5__0_chany_top_out[0:95]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_A1_o_0_(grid_bram_0_right_width_0_height_3_subtile_0__pin_RDATA_A2_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_A1_o_1_(grid_bram_0_right_width_0_height_3_subtile_0__pin_RDATA_A2_o_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_A1_o_2_(grid_bram_0_right_width_0_height_3_subtile_0__pin_RDATA_A2_o_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_A1_o_3_(grid_bram_0_right_width_0_height_3_subtile_0__pin_RDATA_A2_o_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_A1_o_4_(grid_bram_0_right_width_0_height_3_subtile_0__pin_RDATA_A2_o_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_A1_o_5_(grid_bram_0_right_width_0_height_3_subtile_0__pin_RDATA_A2_o_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_B1_o_0_(grid_bram_0_right_width_0_height_3_subtile_0__pin_RDATA_B2_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_B1_o_1_(grid_bram_0_right_width_0_height_3_subtile_0__pin_RDATA_B2_o_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_B1_o_2_(grid_bram_0_right_width_0_height_3_subtile_0__pin_RDATA_B2_o_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_B1_o_3_(grid_bram_0_right_width_0_height_3_subtile_0__pin_RDATA_B2_o_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_B1_o_4_(grid_bram_0_right_width_0_height_3_subtile_0__pin_RDATA_B2_o_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_B1_o_5_(grid_bram_0_right_width_0_height_3_subtile_0__pin_RDATA_B2_o_5_),
		.chanx_left_in(cbx_1__0__27_chanx_right_out[0:95]),
		.ccff_head(grid_clb_28_ccff_tail),
		.chany_top_out(sb_7__2__3_chany_top_out[0:95]),
		.chanx_right_out(sb_7__2__3_chanx_right_out[0:95]),
		.chany_bottom_out(sb_7__2__3_chany_bottom_out[0:95]),
		.chanx_left_out(sb_7__2__3_chanx_left_out[0:95]),
		.ccff_tail(sb_7__2__3_ccff_tail));

	sb_7__2_ sb_7__6_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_7__7__0_chany_bottom_out[0:95]),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_A1_o_6_(grid_bram_0_right_width_0_height_5_subtile_0__pin_RDATA_A2_o_12_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_A1_o_7_(grid_bram_0_right_width_0_height_5_subtile_0__pin_RDATA_A2_o_13_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_A1_o_8_(grid_bram_0_right_width_0_height_5_subtile_0__pin_RDATA_A2_o_14_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_A1_o_9_(grid_bram_0_right_width_0_height_5_subtile_0__pin_RDATA_A2_o_15_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_A1_o_10_(grid_bram_0_right_width_0_height_5_subtile_0__pin_RDATA_A2_o_16_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_A1_o_11_(grid_bram_0_right_width_0_height_5_subtile_0__pin_RDATA_A2_o_17_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_B1_o_6_(grid_bram_0_right_width_0_height_5_subtile_0__pin_RDATA_B2_o_12_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_B1_o_7_(grid_bram_0_right_width_0_height_5_subtile_0__pin_RDATA_B2_o_13_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_B1_o_8_(grid_bram_0_right_width_0_height_5_subtile_0__pin_RDATA_B2_o_14_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_B1_o_9_(grid_bram_0_right_width_0_height_5_subtile_0__pin_RDATA_B2_o_15_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_B1_o_10_(grid_bram_0_right_width_0_height_5_subtile_0__pin_RDATA_B2_o_16_),
		.top_left_grid_right_width_0_height_1_subtile_0__pin_RDATA_B1_o_11_(grid_bram_0_right_width_0_height_5_subtile_0__pin_RDATA_B2_o_17_),
		.chanx_right_in(cbx_2__2__24_chanx_left_out[0:95]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_9_),
		.chany_bottom_in(cby_7__6__0_chany_top_out[0:95]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_A1_o_0_(grid_bram_0_right_width_0_height_4_subtile_0__pin_RDATA_A2_o_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_A1_o_1_(grid_bram_0_right_width_0_height_4_subtile_0__pin_RDATA_A2_o_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_A1_o_2_(grid_bram_0_right_width_0_height_4_subtile_0__pin_RDATA_A2_o_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_A1_o_3_(grid_bram_0_right_width_0_height_4_subtile_0__pin_RDATA_A2_o_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_A1_o_4_(grid_bram_0_right_width_0_height_4_subtile_0__pin_RDATA_A2_o_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_A1_o_5_(grid_bram_0_right_width_0_height_4_subtile_0__pin_RDATA_A2_o_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_B1_o_0_(grid_bram_0_right_width_0_height_4_subtile_0__pin_RDATA_B2_o_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_B1_o_1_(grid_bram_0_right_width_0_height_4_subtile_0__pin_RDATA_B2_o_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_B1_o_2_(grid_bram_0_right_width_0_height_4_subtile_0__pin_RDATA_B2_o_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_B1_o_3_(grid_bram_0_right_width_0_height_4_subtile_0__pin_RDATA_B2_o_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_B1_o_4_(grid_bram_0_right_width_0_height_4_subtile_0__pin_RDATA_B2_o_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_RDATA_B1_o_5_(grid_bram_0_right_width_0_height_4_subtile_0__pin_RDATA_B2_o_11_),
		.chanx_left_in(cbx_1__0__28_chanx_right_out[0:95]),
		.ccff_head(grid_clb_23_ccff_tail),
		.chany_top_out(sb_7__2__4_chany_top_out[0:95]),
		.chanx_right_out(sb_7__2__4_chanx_right_out[0:95]),
		.chany_bottom_out(sb_7__2__4_chany_bottom_out[0:95]),
		.chanx_left_out(sb_7__2__4_chanx_left_out[0:95]),
		.ccff_tail(sb_7__2__4_ccff_tail));

	sb_7__7_ sb_7__7_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_0__1__19_chany_bottom_out[0:95]),
		.chanx_right_in(cbx_2__7__4_chanx_left_out[0:95]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_top_6_bottom_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_9_),
		.chany_bottom_in(cby_7__7__0_chany_top_out[0:95]),
		.bottom_left_grid_right_width_0_height_5_subtile_0__pin_RDATA_A2_o_12_(grid_bram_0_right_width_0_height_5_subtile_0__pin_RDATA_A2_o_12_),
		.bottom_left_grid_right_width_0_height_5_subtile_0__pin_RDATA_A2_o_13_(grid_bram_0_right_width_0_height_5_subtile_0__pin_RDATA_A2_o_13_),
		.bottom_left_grid_right_width_0_height_5_subtile_0__pin_RDATA_A2_o_14_(grid_bram_0_right_width_0_height_5_subtile_0__pin_RDATA_A2_o_14_),
		.bottom_left_grid_right_width_0_height_5_subtile_0__pin_RDATA_A2_o_15_(grid_bram_0_right_width_0_height_5_subtile_0__pin_RDATA_A2_o_15_),
		.bottom_left_grid_right_width_0_height_5_subtile_0__pin_RDATA_A2_o_16_(grid_bram_0_right_width_0_height_5_subtile_0__pin_RDATA_A2_o_16_),
		.bottom_left_grid_right_width_0_height_5_subtile_0__pin_RDATA_A2_o_17_(grid_bram_0_right_width_0_height_5_subtile_0__pin_RDATA_A2_o_17_),
		.bottom_left_grid_right_width_0_height_5_subtile_0__pin_RDATA_B2_o_12_(grid_bram_0_right_width_0_height_5_subtile_0__pin_RDATA_B2_o_12_),
		.bottom_left_grid_right_width_0_height_5_subtile_0__pin_RDATA_B2_o_13_(grid_bram_0_right_width_0_height_5_subtile_0__pin_RDATA_B2_o_13_),
		.bottom_left_grid_right_width_0_height_5_subtile_0__pin_RDATA_B2_o_14_(grid_bram_0_right_width_0_height_5_subtile_0__pin_RDATA_B2_o_14_),
		.bottom_left_grid_right_width_0_height_5_subtile_0__pin_RDATA_B2_o_15_(grid_bram_0_right_width_0_height_5_subtile_0__pin_RDATA_B2_o_15_),
		.bottom_left_grid_right_width_0_height_5_subtile_0__pin_RDATA_B2_o_16_(grid_bram_0_right_width_0_height_5_subtile_0__pin_RDATA_B2_o_16_),
		.bottom_left_grid_right_width_0_height_5_subtile_0__pin_RDATA_B2_o_17_(grid_bram_0_right_width_0_height_5_subtile_0__pin_RDATA_B2_o_17_),
		.chanx_left_in(cbx_4__7__1_chanx_right_out[0:95]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_top_5_bottom_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.ccff_head(grid_io_top_6_ccff_tail),
		.chany_top_out(sb_7__7__0_chany_top_out[0:95]),
		.chanx_right_out(sb_7__7__0_chanx_right_out[0:95]),
		.chany_bottom_out(sb_7__7__0_chany_bottom_out[0:95]),
		.chanx_left_out(sb_7__7__0_chanx_left_out[0:95]),
		.ccff_tail(sb_7__7__0_ccff_tail));

	sb_9__1_ sb_9__1_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_9__2__0_chany_bottom_out[0:95]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_16_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_18_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_19_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.chanx_right_in(cbx_1__0__35_chanx_left_out[0:95]),
		.chany_bottom_in(cby_9__1__0_chany_top_out[0:95]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_right_0_left_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.chanx_left_in(cbx_2__1__5_chanx_right_out[0:95]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_bottom_7_top_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.ccff_head(grid_io_right_1_ccff_tail),
		.chany_top_out(sb_9__1__0_chany_top_out[0:95]),
		.chanx_right_out(sb_9__1__0_chanx_right_out[0:95]),
		.chany_bottom_out(sb_9__1__0_chany_bottom_out[0:95]),
		.chanx_left_out(sb_9__1__0_chanx_left_out[0:95]),
		.ccff_tail(sb_9__1__0_ccff_tail));

	sb_9__2_ sb_9__2_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_9__2__1_chany_bottom_out[0:95]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_16_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_18_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_19_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.chanx_right_in(cbx_1__0__36_chanx_left_out[0:95]),
		.chany_bottom_in(cby_9__2__0_chany_top_out[0:95]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_right_1_left_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_left_in(cbx_2__2__25_chanx_right_out[0:95]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_7_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_9_),
		.ccff_head(grid_clb_25_ccff_tail),
		.chany_top_out(sb_9__2__0_chany_top_out[0:95]),
		.chanx_right_out(sb_9__2__0_chanx_right_out[0:95]),
		.chany_bottom_out(sb_9__2__0_chany_bottom_out[0:95]),
		.chanx_left_out(sb_9__2__0_chanx_left_out[0:95]),
		.ccff_tail(sb_9__2__0_ccff_tail));

	sb_9__2_ sb_9__3_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_9__2__2_chany_bottom_out[0:95]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_16_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_18_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_19_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.chanx_right_in(cbx_1__0__37_chanx_left_out[0:95]),
		.chany_bottom_in(cby_9__2__1_chany_top_out[0:95]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_right_2_left_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_left_in(cbx_2__2__26_chanx_right_out[0:95]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_7_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_9_),
		.ccff_head(grid_io_right_3_ccff_tail),
		.chany_top_out(sb_9__2__1_chany_top_out[0:95]),
		.chanx_right_out(sb_9__2__1_chanx_right_out[0:95]),
		.chany_bottom_out(sb_9__2__1_chany_bottom_out[0:95]),
		.chanx_left_out(sb_9__2__1_chanx_left_out[0:95]),
		.ccff_tail(sb_9__2__1_ccff_tail));

	sb_9__2_ sb_9__4_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_9__2__3_chany_bottom_out[0:95]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_16_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_18_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_19_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.chanx_right_in(cbx_1__0__38_chanx_left_out[0:95]),
		.chany_bottom_in(cby_9__2__2_chany_top_out[0:95]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_right_3_left_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_left_in(cbx_2__2__27_chanx_right_out[0:95]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_7_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_9_),
		.ccff_head(grid_clb_27_ccff_tail),
		.chany_top_out(sb_9__2__2_chany_top_out[0:95]),
		.chanx_right_out(sb_9__2__2_chanx_right_out[0:95]),
		.chany_bottom_out(sb_9__2__2_chany_bottom_out[0:95]),
		.chanx_left_out(sb_9__2__2_chanx_left_out[0:95]),
		.ccff_tail(sb_9__2__2_ccff_tail));

	sb_9__2_ sb_9__5_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_9__2__4_chany_bottom_out[0:95]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_16_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_18_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_19_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.chanx_right_in(cbx_1__0__39_chanx_left_out[0:95]),
		.chany_bottom_in(cby_9__2__3_chany_top_out[0:95]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_right_4_left_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_left_in(cbx_2__2__28_chanx_right_out[0:95]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_7_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_9_),
		.ccff_head(grid_io_right_5_ccff_tail),
		.chany_top_out(sb_9__2__3_chany_top_out[0:95]),
		.chanx_right_out(sb_9__2__3_chanx_right_out[0:95]),
		.chany_bottom_out(sb_9__2__3_chany_bottom_out[0:95]),
		.chanx_left_out(sb_9__2__3_chanx_left_out[0:95]),
		.ccff_tail(sb_9__2__3_ccff_tail));

	sb_9__2_ sb_9__6_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_9__2__5_chany_bottom_out[0:95]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_16_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_17_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_18_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_19_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.chanx_right_in(cbx_1__0__40_chanx_left_out[0:95]),
		.chany_bottom_in(cby_9__2__4_chany_top_out[0:95]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_right_5_left_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_left_in(cbx_2__2__29_chanx_right_out[0:95]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_7_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_9_),
		.ccff_head(grid_clb_29_ccff_tail),
		.chany_top_out(sb_9__2__4_chany_top_out[0:95]),
		.chanx_right_out(sb_9__2__4_chanx_right_out[0:95]),
		.chany_bottom_out(sb_9__2__4_chany_bottom_out[0:95]),
		.chanx_left_out(sb_9__2__4_chanx_left_out[0:95]),
		.ccff_tail(sb_9__2__4_ccff_tail));

	sb_9__7_ sb_9__7_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_9__1__1_chany_bottom_out[0:95]),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.top_right_grid_left_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_right_7_left_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.chanx_right_in(cbx_1__0__41_chanx_left_out[0:95]),
		.chany_bottom_in(cby_9__2__5_chany_top_out[0:95]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_right_6_left_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_16_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_17_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_18_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_19_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_19_),
		.chanx_left_in(cbx_2__7__5_chanx_right_out[0:95]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_8__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_8__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_9__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_9__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_10__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_10__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_11__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_11__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_12__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_12__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_13__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_13__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_14__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_14__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_15__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_15__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_16__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_16__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_17__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_17__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_18__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_18__pin_a2f_o_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_19__pin_a2f_o_0_(grid_io_top_7_bottom_width_0_height_0_subtile_19__pin_a2f_o_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_7_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_9_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_9_),
		.ccff_head(ccff_head[9]),
		.chany_top_out(sb_9__7__0_chany_top_out[0:95]),
		.chanx_right_out(sb_9__7__0_chanx_right_out[0:95]),
		.chany_bottom_out(sb_9__7__0_chany_bottom_out[0:95]),
		.chanx_left_out(sb_9__7__0_chanx_left_out[0:95]),
		.ccff_tail(sb_9__7__0_ccff_tail));

	sb_10__0_ sb_10__0_ (
		.chany_top_in(cby_0__1__22_chany_bottom_out[0:95]),
		.chanx_left_in(cbx_1__0__34_chanx_right_out[0:95]),
		.chany_top_out(sb_10__0__0_chany_top_out[0:95]),
		.chanx_left_out(sb_10__0__0_chanx_left_out[0:95]));

	sb_10__1_ sb_10__1_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_0__1__23_chany_bottom_out[0:95]),
		.chany_bottom_in(cby_0__1__22_chany_top_out[0:95]),
		.chanx_left_in(cbx_1__0__35_chanx_right_out[0:95]),
		.ccff_head(grid_io_right_0_ccff_tail),
		.chany_top_out(sb_10__1__0_chany_top_out[0:95]),
		.chany_bottom_out(sb_10__1__0_chany_bottom_out[0:95]),
		.chanx_left_out(sb_10__1__0_chanx_left_out[0:95]),
		.ccff_tail(sb_10__1__0_ccff_tail));

	sb_10__1_ sb_10__2_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_0__1__24_chany_bottom_out[0:95]),
		.chany_bottom_in(cby_0__1__23_chany_top_out[0:95]),
		.chanx_left_in(cbx_1__0__36_chanx_right_out[0:95]),
		.ccff_head(grid_clb_31_ccff_tail),
		.chany_top_out(sb_10__1__1_chany_top_out[0:95]),
		.chany_bottom_out(sb_10__1__1_chany_bottom_out[0:95]),
		.chanx_left_out(sb_10__1__1_chanx_left_out[0:95]),
		.ccff_tail(sb_10__1__1_ccff_tail));

	sb_10__1_ sb_10__3_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_0__1__25_chany_bottom_out[0:95]),
		.chany_bottom_in(cby_0__1__24_chany_top_out[0:95]),
		.chanx_left_in(cbx_1__0__37_chanx_right_out[0:95]),
		.ccff_head(grid_io_right_2_ccff_tail),
		.chany_top_out(sb_10__1__2_chany_top_out[0:95]),
		.chany_bottom_out(sb_10__1__2_chany_bottom_out[0:95]),
		.chanx_left_out(sb_10__1__2_chanx_left_out[0:95]),
		.ccff_tail(ccff_tail[3]));

	sb_10__1_ sb_10__4_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_0__1__26_chany_bottom_out[0:95]),
		.chany_bottom_in(cby_0__1__25_chany_top_out[0:95]),
		.chanx_left_in(cbx_1__0__38_chanx_right_out[0:95]),
		.ccff_head(grid_clb_33_ccff_tail),
		.chany_top_out(sb_10__1__3_chany_top_out[0:95]),
		.chany_bottom_out(sb_10__1__3_chany_bottom_out[0:95]),
		.chanx_left_out(sb_10__1__3_chanx_left_out[0:95]),
		.ccff_tail(sb_10__1__3_ccff_tail));

	sb_10__1_ sb_10__5_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_0__1__27_chany_bottom_out[0:95]),
		.chany_bottom_in(cby_0__1__26_chany_top_out[0:95]),
		.chanx_left_in(cbx_1__0__39_chanx_right_out[0:95]),
		.ccff_head(grid_io_right_4_ccff_tail),
		.chany_top_out(sb_10__1__4_chany_top_out[0:95]),
		.chany_bottom_out(sb_10__1__4_chany_bottom_out[0:95]),
		.chanx_left_out(sb_10__1__4_chanx_left_out[0:95]),
		.ccff_tail(sb_10__1__4_ccff_tail));

	sb_10__1_ sb_10__6_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_0__1__28_chany_bottom_out[0:95]),
		.chany_bottom_in(cby_0__1__27_chany_top_out[0:95]),
		.chanx_left_in(cbx_1__0__40_chanx_right_out[0:95]),
		.ccff_head(grid_clb_35_ccff_tail),
		.chany_top_out(sb_10__1__5_chany_top_out[0:95]),
		.chany_bottom_out(sb_10__1__5_chany_bottom_out[0:95]),
		.chanx_left_out(sb_10__1__5_chanx_left_out[0:95]),
		.ccff_tail(sb_10__1__5_ccff_tail));

	sb_10__1_ sb_10__7_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_top_in(cby_0__1__29_chany_bottom_out[0:95]),
		.chany_bottom_in(cby_0__1__28_chany_top_out[0:95]),
		.chanx_left_in(cbx_1__0__41_chanx_right_out[0:95]),
		.ccff_head(grid_io_right_6_ccff_tail),
		.chany_top_out(sb_10__1__6_chany_top_out[0:95]),
		.chany_bottom_out(sb_10__1__6_chany_bottom_out[0:95]),
		.chanx_left_out(sb_10__1__6_chanx_left_out[0:95]),
		.ccff_tail(sb_10__1__6_ccff_tail));

	sb_10__8_ sb_10__8_ (
		.chany_bottom_in(cby_0__1__29_chany_top_out[0:95]),
		.chanx_left_in(cbx_1__0__42_chanx_right_out[0:95]),
		.chany_bottom_out(sb_10__8__0_chany_bottom_out[0:95]),
		.chanx_left_out(sb_10__8__0_chanx_left_out[0:95]));

	cbx_1__0_ cbx_1__0_ (
		.chanx_left_in(sb_0__0__0_chanx_right_out[0:95]),
		.chanx_right_in(sb_1__0__0_chanx_left_out[0:95]),
		.chanx_left_out(cbx_1__0__0_chanx_left_out[0:95]),
		.chanx_right_out(cbx_1__0__0_chanx_right_out[0:95]));

	cbx_1__0_ cbx_1__1_ (
		.chanx_left_in(sb_0__1__0_chanx_right_out[0:95]),
		.chanx_right_in(sb_1__1__0_chanx_left_out[0:95]),
		.chanx_left_out(cbx_1__0__1_chanx_left_out[0:95]),
		.chanx_right_out(cbx_1__0__1_chanx_right_out[0:95]));

	cbx_1__0_ cbx_1__2_ (
		.chanx_left_in(sb_0__1__1_chanx_right_out[0:95]),
		.chanx_right_in(sb_1__2__0_chanx_left_out[0:95]),
		.chanx_left_out(cbx_1__0__2_chanx_left_out[0:95]),
		.chanx_right_out(cbx_1__0__2_chanx_right_out[0:95]));

	cbx_1__0_ cbx_1__3_ (
		.chanx_left_in(sb_0__1__2_chanx_right_out[0:95]),
		.chanx_right_in(sb_1__2__1_chanx_left_out[0:95]),
		.chanx_left_out(cbx_1__0__3_chanx_left_out[0:95]),
		.chanx_right_out(cbx_1__0__3_chanx_right_out[0:95]));

	cbx_1__0_ cbx_1__4_ (
		.chanx_left_in(sb_0__1__3_chanx_right_out[0:95]),
		.chanx_right_in(sb_1__2__2_chanx_left_out[0:95]),
		.chanx_left_out(cbx_1__0__4_chanx_left_out[0:95]),
		.chanx_right_out(cbx_1__0__4_chanx_right_out[0:95]));

	cbx_1__0_ cbx_1__5_ (
		.chanx_left_in(sb_0__1__4_chanx_right_out[0:95]),
		.chanx_right_in(sb_1__2__3_chanx_left_out[0:95]),
		.chanx_left_out(cbx_1__0__5_chanx_left_out[0:95]),
		.chanx_right_out(cbx_1__0__5_chanx_right_out[0:95]));

	cbx_1__0_ cbx_1__6_ (
		.chanx_left_in(sb_0__1__5_chanx_right_out[0:95]),
		.chanx_right_in(sb_1__2__4_chanx_left_out[0:95]),
		.chanx_left_out(cbx_1__0__6_chanx_left_out[0:95]),
		.chanx_right_out(cbx_1__0__6_chanx_right_out[0:95]));

	cbx_1__0_ cbx_1__7_ (
		.chanx_left_in(sb_0__1__6_chanx_right_out[0:95]),
		.chanx_right_in(sb_1__7__0_chanx_left_out[0:95]),
		.chanx_left_out(cbx_1__0__7_chanx_left_out[0:95]),
		.chanx_right_out(cbx_1__0__7_chanx_right_out[0:95]));

	cbx_1__0_ cbx_1__8_ (
		.chanx_left_in(sb_0__8__0_chanx_right_out[0:95]),
		.chanx_right_in(sb_1__8__0_chanx_left_out[0:95]),
		.chanx_left_out(cbx_1__0__8_chanx_left_out[0:95]),
		.chanx_right_out(cbx_1__0__8_chanx_right_out[0:95]));

	cbx_1__0_ cbx_2__0_ (
		.chanx_left_in(sb_1__0__0_chanx_right_out[0:95]),
		.chanx_right_in(sb_2__0__0_chanx_left_out[0:95]),
		.chanx_left_out(cbx_1__0__9_chanx_left_out[0:95]),
		.chanx_right_out(cbx_1__0__9_chanx_right_out[0:95]));

	cbx_1__0_ cbx_2__8_ (
		.chanx_left_in(sb_1__8__0_chanx_right_out[0:95]),
		.chanx_right_in(sb_2__8__0_chanx_left_out[0:95]),
		.chanx_left_out(cbx_1__0__10_chanx_left_out[0:95]),
		.chanx_right_out(cbx_1__0__10_chanx_right_out[0:95]));

	cbx_1__0_ cbx_3__0_ (
		.chanx_left_in(sb_2__0__0_chanx_right_out[0:95]),
		.chanx_right_in(sb_2__0__1_chanx_left_out[0:95]),
		.chanx_left_out(cbx_1__0__11_chanx_left_out[0:95]),
		.chanx_right_out(cbx_1__0__11_chanx_right_out[0:95]));

	cbx_1__0_ cbx_3__8_ (
		.chanx_left_in(sb_2__8__0_chanx_right_out[0:95]),
		.chanx_right_in(sb_2__8__1_chanx_left_out[0:95]),
		.chanx_left_out(cbx_1__0__12_chanx_left_out[0:95]),
		.chanx_right_out(cbx_1__0__12_chanx_right_out[0:95]));

	cbx_1__0_ cbx_4__0_ (
		.chanx_left_in(sb_2__0__1_chanx_right_out[0:95]),
		.chanx_right_in(sb_2__0__2_chanx_left_out[0:95]),
		.chanx_left_out(cbx_1__0__13_chanx_left_out[0:95]),
		.chanx_right_out(cbx_1__0__13_chanx_right_out[0:95]));

	cbx_1__0_ cbx_4__2_ (
		.chanx_left_in(sb_3__2__0_chanx_right_out[0:95]),
		.chanx_right_in(sb_4__2__0_chanx_left_out[0:95]),
		.chanx_left_out(cbx_1__0__14_chanx_left_out[0:95]),
		.chanx_right_out(cbx_1__0__14_chanx_right_out[0:95]));

	cbx_1__0_ cbx_4__3_ (
		.chanx_left_in(sb_3__2__1_chanx_right_out[0:95]),
		.chanx_right_in(sb_4__3__0_chanx_left_out[0:95]),
		.chanx_left_out(cbx_1__0__15_chanx_left_out[0:95]),
		.chanx_right_out(cbx_1__0__15_chanx_right_out[0:95]));

	cbx_1__0_ cbx_4__5_ (
		.chanx_left_in(sb_3__2__2_chanx_right_out[0:95]),
		.chanx_right_in(sb_4__2__1_chanx_left_out[0:95]),
		.chanx_left_out(cbx_1__0__16_chanx_left_out[0:95]),
		.chanx_right_out(cbx_1__0__16_chanx_right_out[0:95]));

	cbx_1__0_ cbx_4__6_ (
		.chanx_left_in(sb_3__2__3_chanx_right_out[0:95]),
		.chanx_right_in(sb_4__3__1_chanx_left_out[0:95]),
		.chanx_left_out(cbx_1__0__17_chanx_left_out[0:95]),
		.chanx_right_out(cbx_1__0__17_chanx_right_out[0:95]));

	cbx_1__0_ cbx_4__8_ (
		.chanx_left_in(sb_2__8__1_chanx_right_out[0:95]),
		.chanx_right_in(sb_2__8__2_chanx_left_out[0:95]),
		.chanx_left_out(cbx_1__0__18_chanx_left_out[0:95]),
		.chanx_right_out(cbx_1__0__18_chanx_right_out[0:95]));

	cbx_1__0_ cbx_5__0_ (
		.chanx_left_in(sb_2__0__2_chanx_right_out[0:95]),
		.chanx_right_in(sb_2__0__3_chanx_left_out[0:95]),
		.chanx_left_out(cbx_1__0__19_chanx_left_out[0:95]),
		.chanx_right_out(cbx_1__0__19_chanx_right_out[0:95]));

	cbx_1__0_ cbx_5__8_ (
		.chanx_left_in(sb_2__8__2_chanx_right_out[0:95]),
		.chanx_right_in(sb_2__8__3_chanx_left_out[0:95]),
		.chanx_left_out(cbx_1__0__20_chanx_left_out[0:95]),
		.chanx_right_out(cbx_1__0__20_chanx_right_out[0:95]));

	cbx_1__0_ cbx_6__0_ (
		.chanx_left_in(sb_2__0__3_chanx_right_out[0:95]),
		.chanx_right_in(sb_2__0__4_chanx_left_out[0:95]),
		.chanx_left_out(cbx_1__0__21_chanx_left_out[0:95]),
		.chanx_right_out(cbx_1__0__21_chanx_right_out[0:95]));

	cbx_1__0_ cbx_6__8_ (
		.chanx_left_in(sb_2__8__3_chanx_right_out[0:95]),
		.chanx_right_in(sb_2__8__4_chanx_left_out[0:95]),
		.chanx_left_out(cbx_1__0__22_chanx_left_out[0:95]),
		.chanx_right_out(cbx_1__0__22_chanx_right_out[0:95]));

	cbx_1__0_ cbx_7__0_ (
		.chanx_left_in(sb_2__0__4_chanx_right_out[0:95]),
		.chanx_right_in(sb_2__0__5_chanx_left_out[0:95]),
		.chanx_left_out(cbx_1__0__23_chanx_left_out[0:95]),
		.chanx_right_out(cbx_1__0__23_chanx_right_out[0:95]));

	cbx_1__0_ cbx_7__2_ (
		.chanx_left_in(sb_3__2__4_chanx_right_out[0:95]),
		.chanx_right_in(sb_7__2__0_chanx_left_out[0:95]),
		.chanx_left_out(cbx_1__0__24_chanx_left_out[0:95]),
		.chanx_right_out(cbx_1__0__24_chanx_right_out[0:95]));

	cbx_1__0_ cbx_7__3_ (
		.chanx_left_in(sb_3__2__5_chanx_right_out[0:95]),
		.chanx_right_in(sb_7__2__1_chanx_left_out[0:95]),
		.chanx_left_out(cbx_1__0__25_chanx_left_out[0:95]),
		.chanx_right_out(cbx_1__0__25_chanx_right_out[0:95]));

	cbx_1__0_ cbx_7__4_ (
		.chanx_left_in(sb_3__2__6_chanx_right_out[0:95]),
		.chanx_right_in(sb_7__2__2_chanx_left_out[0:95]),
		.chanx_left_out(cbx_1__0__26_chanx_left_out[0:95]),
		.chanx_right_out(cbx_1__0__26_chanx_right_out[0:95]));

	cbx_1__0_ cbx_7__5_ (
		.chanx_left_in(sb_3__2__7_chanx_right_out[0:95]),
		.chanx_right_in(sb_7__2__3_chanx_left_out[0:95]),
		.chanx_left_out(cbx_1__0__27_chanx_left_out[0:95]),
		.chanx_right_out(cbx_1__0__27_chanx_right_out[0:95]));

	cbx_1__0_ cbx_7__6_ (
		.chanx_left_in(sb_3__2__8_chanx_right_out[0:95]),
		.chanx_right_in(sb_7__2__4_chanx_left_out[0:95]),
		.chanx_left_out(cbx_1__0__28_chanx_left_out[0:95]),
		.chanx_right_out(cbx_1__0__28_chanx_right_out[0:95]));

	cbx_1__0_ cbx_7__8_ (
		.chanx_left_in(sb_2__8__4_chanx_right_out[0:95]),
		.chanx_right_in(sb_2__8__5_chanx_left_out[0:95]),
		.chanx_left_out(cbx_1__0__29_chanx_left_out[0:95]),
		.chanx_right_out(cbx_1__0__29_chanx_right_out[0:95]));

	cbx_1__0_ cbx_8__0_ (
		.chanx_left_in(sb_2__0__5_chanx_right_out[0:95]),
		.chanx_right_in(sb_2__0__6_chanx_left_out[0:95]),
		.chanx_left_out(cbx_1__0__30_chanx_left_out[0:95]),
		.chanx_right_out(cbx_1__0__30_chanx_right_out[0:95]));

	cbx_1__0_ cbx_8__8_ (
		.chanx_left_in(sb_2__8__5_chanx_right_out[0:95]),
		.chanx_right_in(sb_2__8__6_chanx_left_out[0:95]),
		.chanx_left_out(cbx_1__0__31_chanx_left_out[0:95]),
		.chanx_right_out(cbx_1__0__31_chanx_right_out[0:95]));

	cbx_1__0_ cbx_9__0_ (
		.chanx_left_in(sb_2__0__6_chanx_right_out[0:95]),
		.chanx_right_in(sb_1__0__1_chanx_left_out[0:95]),
		.chanx_left_out(cbx_1__0__32_chanx_left_out[0:95]),
		.chanx_right_out(cbx_1__0__32_chanx_right_out[0:95]));

	cbx_1__0_ cbx_9__8_ (
		.chanx_left_in(sb_2__8__6_chanx_right_out[0:95]),
		.chanx_right_in(sb_1__8__1_chanx_left_out[0:95]),
		.chanx_left_out(cbx_1__0__33_chanx_left_out[0:95]),
		.chanx_right_out(cbx_1__0__33_chanx_right_out[0:95]));

	cbx_1__0_ cbx_10__0_ (
		.chanx_left_in(sb_1__0__1_chanx_right_out[0:95]),
		.chanx_right_in(sb_10__0__0_chanx_left_out[0:95]),
		.chanx_left_out(cbx_1__0__34_chanx_left_out[0:95]),
		.chanx_right_out(cbx_1__0__34_chanx_right_out[0:95]));

	cbx_1__0_ cbx_10__1_ (
		.chanx_left_in(sb_9__1__0_chanx_right_out[0:95]),
		.chanx_right_in(sb_10__1__0_chanx_left_out[0:95]),
		.chanx_left_out(cbx_1__0__35_chanx_left_out[0:95]),
		.chanx_right_out(cbx_1__0__35_chanx_right_out[0:95]));

	cbx_1__0_ cbx_10__2_ (
		.chanx_left_in(sb_9__2__0_chanx_right_out[0:95]),
		.chanx_right_in(sb_10__1__1_chanx_left_out[0:95]),
		.chanx_left_out(cbx_1__0__36_chanx_left_out[0:95]),
		.chanx_right_out(cbx_1__0__36_chanx_right_out[0:95]));

	cbx_1__0_ cbx_10__3_ (
		.chanx_left_in(sb_9__2__1_chanx_right_out[0:95]),
		.chanx_right_in(sb_10__1__2_chanx_left_out[0:95]),
		.chanx_left_out(cbx_1__0__37_chanx_left_out[0:95]),
		.chanx_right_out(cbx_1__0__37_chanx_right_out[0:95]));

	cbx_1__0_ cbx_10__4_ (
		.chanx_left_in(sb_9__2__2_chanx_right_out[0:95]),
		.chanx_right_in(sb_10__1__3_chanx_left_out[0:95]),
		.chanx_left_out(cbx_1__0__38_chanx_left_out[0:95]),
		.chanx_right_out(cbx_1__0__38_chanx_right_out[0:95]));

	cbx_1__0_ cbx_10__5_ (
		.chanx_left_in(sb_9__2__3_chanx_right_out[0:95]),
		.chanx_right_in(sb_10__1__4_chanx_left_out[0:95]),
		.chanx_left_out(cbx_1__0__39_chanx_left_out[0:95]),
		.chanx_right_out(cbx_1__0__39_chanx_right_out[0:95]));

	cbx_1__0_ cbx_10__6_ (
		.chanx_left_in(sb_9__2__4_chanx_right_out[0:95]),
		.chanx_right_in(sb_10__1__5_chanx_left_out[0:95]),
		.chanx_left_out(cbx_1__0__40_chanx_left_out[0:95]),
		.chanx_right_out(cbx_1__0__40_chanx_right_out[0:95]));

	cbx_1__0_ cbx_10__7_ (
		.chanx_left_in(sb_9__7__0_chanx_right_out[0:95]),
		.chanx_right_in(sb_10__1__6_chanx_left_out[0:95]),
		.chanx_left_out(cbx_1__0__41_chanx_left_out[0:95]),
		.chanx_right_out(cbx_1__0__41_chanx_right_out[0:95]));

	cbx_1__0_ cbx_10__8_ (
		.chanx_left_in(sb_1__8__1_chanx_right_out[0:95]),
		.chanx_right_in(sb_10__8__0_chanx_left_out[0:95]),
		.chanx_left_out(cbx_1__0__42_chanx_left_out[0:95]),
		.chanx_right_out(cbx_1__0__42_chanx_right_out[0:95]));

	cbx_2__1_ cbx_2__1_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chanx_left_in(sb_1__1__0_chanx_right_out[0:95]),
		.chanx_right_in(sb_2__1__0_chanx_left_out[0:95]),
		.ccff_head(sb_2__1__0_ccff_tail),
		.chanx_left_out(cbx_2__1__0_chanx_left_out[0:95]),
		.chanx_right_out(cbx_2__1__0_chanx_right_out[0:95]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_f2a_i_0_(cbx_2__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_f2a_i_0_(cbx_2__1__0_bottom_grid_top_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_f2a_i_0_(cbx_2__1__0_bottom_grid_top_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_f2a_i_0_(cbx_2__1__0_bottom_grid_top_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_f2a_i_0_(cbx_2__1__0_bottom_grid_top_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_f2a_i_0_(cbx_2__1__0_bottom_grid_top_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_f2a_i_0_(cbx_2__1__0_bottom_grid_top_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_f2a_i_0_(cbx_2__1__0_bottom_grid_top_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_f2a_i_0_(cbx_2__1__0_bottom_grid_top_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_9__pin_f2a_i_0_(cbx_2__1__0_bottom_grid_top_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_10__pin_f2a_i_0_(cbx_2__1__0_bottom_grid_top_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_11__pin_f2a_i_0_(cbx_2__1__0_bottom_grid_top_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_12__pin_f2a_i_0_(cbx_2__1__0_bottom_grid_top_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_13__pin_f2a_i_0_(cbx_2__1__0_bottom_grid_top_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_14__pin_f2a_i_0_(cbx_2__1__0_bottom_grid_top_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_15__pin_f2a_i_0_(cbx_2__1__0_bottom_grid_top_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_16__pin_f2a_i_0_(cbx_2__1__0_bottom_grid_top_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_17__pin_f2a_i_0_(cbx_2__1__0_bottom_grid_top_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_18__pin_f2a_i_0_(cbx_2__1__0_bottom_grid_top_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_19__pin_f2a_i_0_(cbx_2__1__0_bottom_grid_top_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.ccff_tail(cbx_2__1__0_ccff_tail));

	cbx_2__1_ cbx_3__1_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chanx_left_in(sb_2__1__0_chanx_right_out[0:95]),
		.chanx_right_in(sb_3__1__0_chanx_left_out[0:95]),
		.ccff_head(sb_3__1__0_ccff_tail),
		.chanx_left_out(cbx_2__1__1_chanx_left_out[0:95]),
		.chanx_right_out(cbx_2__1__1_chanx_right_out[0:95]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_f2a_i_0_(cbx_2__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_f2a_i_0_(cbx_2__1__1_bottom_grid_top_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_f2a_i_0_(cbx_2__1__1_bottom_grid_top_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_f2a_i_0_(cbx_2__1__1_bottom_grid_top_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_f2a_i_0_(cbx_2__1__1_bottom_grid_top_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_f2a_i_0_(cbx_2__1__1_bottom_grid_top_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_f2a_i_0_(cbx_2__1__1_bottom_grid_top_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_f2a_i_0_(cbx_2__1__1_bottom_grid_top_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_f2a_i_0_(cbx_2__1__1_bottom_grid_top_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_9__pin_f2a_i_0_(cbx_2__1__1_bottom_grid_top_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_10__pin_f2a_i_0_(cbx_2__1__1_bottom_grid_top_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_11__pin_f2a_i_0_(cbx_2__1__1_bottom_grid_top_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_12__pin_f2a_i_0_(cbx_2__1__1_bottom_grid_top_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_13__pin_f2a_i_0_(cbx_2__1__1_bottom_grid_top_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_14__pin_f2a_i_0_(cbx_2__1__1_bottom_grid_top_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_15__pin_f2a_i_0_(cbx_2__1__1_bottom_grid_top_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_16__pin_f2a_i_0_(cbx_2__1__1_bottom_grid_top_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_17__pin_f2a_i_0_(cbx_2__1__1_bottom_grid_top_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_18__pin_f2a_i_0_(cbx_2__1__1_bottom_grid_top_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_19__pin_f2a_i_0_(cbx_2__1__1_bottom_grid_top_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.ccff_tail(cbx_2__1__1_ccff_tail));

	cbx_2__1_ cbx_5__1_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chanx_left_in(sb_4__1__0_chanx_right_out[0:95]),
		.chanx_right_in(sb_2__1__1_chanx_left_out[0:95]),
		.ccff_head(sb_2__1__1_ccff_tail),
		.chanx_left_out(cbx_2__1__2_chanx_left_out[0:95]),
		.chanx_right_out(cbx_2__1__2_chanx_right_out[0:95]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_f2a_i_0_(cbx_2__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_f2a_i_0_(cbx_2__1__2_bottom_grid_top_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_f2a_i_0_(cbx_2__1__2_bottom_grid_top_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_f2a_i_0_(cbx_2__1__2_bottom_grid_top_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_f2a_i_0_(cbx_2__1__2_bottom_grid_top_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_f2a_i_0_(cbx_2__1__2_bottom_grid_top_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_f2a_i_0_(cbx_2__1__2_bottom_grid_top_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_f2a_i_0_(cbx_2__1__2_bottom_grid_top_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_f2a_i_0_(cbx_2__1__2_bottom_grid_top_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_9__pin_f2a_i_0_(cbx_2__1__2_bottom_grid_top_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_10__pin_f2a_i_0_(cbx_2__1__2_bottom_grid_top_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_11__pin_f2a_i_0_(cbx_2__1__2_bottom_grid_top_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_12__pin_f2a_i_0_(cbx_2__1__2_bottom_grid_top_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_13__pin_f2a_i_0_(cbx_2__1__2_bottom_grid_top_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_14__pin_f2a_i_0_(cbx_2__1__2_bottom_grid_top_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_15__pin_f2a_i_0_(cbx_2__1__2_bottom_grid_top_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_16__pin_f2a_i_0_(cbx_2__1__2_bottom_grid_top_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_17__pin_f2a_i_0_(cbx_2__1__2_bottom_grid_top_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_18__pin_f2a_i_0_(cbx_2__1__2_bottom_grid_top_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_19__pin_f2a_i_0_(cbx_2__1__2_bottom_grid_top_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.ccff_tail(cbx_2__1__2_ccff_tail));

	cbx_2__1_ cbx_6__1_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chanx_left_in(sb_2__1__1_chanx_right_out[0:95]),
		.chanx_right_in(sb_2__1__2_chanx_left_out[0:95]),
		.ccff_head(sb_2__1__2_ccff_tail),
		.chanx_left_out(cbx_2__1__3_chanx_left_out[0:95]),
		.chanx_right_out(cbx_2__1__3_chanx_right_out[0:95]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_f2a_i_0_(cbx_2__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_f2a_i_0_(cbx_2__1__3_bottom_grid_top_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_f2a_i_0_(cbx_2__1__3_bottom_grid_top_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_f2a_i_0_(cbx_2__1__3_bottom_grid_top_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_f2a_i_0_(cbx_2__1__3_bottom_grid_top_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_f2a_i_0_(cbx_2__1__3_bottom_grid_top_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_f2a_i_0_(cbx_2__1__3_bottom_grid_top_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_f2a_i_0_(cbx_2__1__3_bottom_grid_top_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_f2a_i_0_(cbx_2__1__3_bottom_grid_top_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_9__pin_f2a_i_0_(cbx_2__1__3_bottom_grid_top_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_10__pin_f2a_i_0_(cbx_2__1__3_bottom_grid_top_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_11__pin_f2a_i_0_(cbx_2__1__3_bottom_grid_top_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_12__pin_f2a_i_0_(cbx_2__1__3_bottom_grid_top_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_13__pin_f2a_i_0_(cbx_2__1__3_bottom_grid_top_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_14__pin_f2a_i_0_(cbx_2__1__3_bottom_grid_top_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_15__pin_f2a_i_0_(cbx_2__1__3_bottom_grid_top_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_16__pin_f2a_i_0_(cbx_2__1__3_bottom_grid_top_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_17__pin_f2a_i_0_(cbx_2__1__3_bottom_grid_top_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_18__pin_f2a_i_0_(cbx_2__1__3_bottom_grid_top_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_19__pin_f2a_i_0_(cbx_2__1__3_bottom_grid_top_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.ccff_tail(cbx_2__1__3_ccff_tail));

	cbx_2__1_ cbx_8__1_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chanx_left_in(sb_7__1__0_chanx_right_out[0:95]),
		.chanx_right_in(sb_2__1__3_chanx_left_out[0:95]),
		.ccff_head(sb_2__1__3_ccff_tail),
		.chanx_left_out(cbx_2__1__4_chanx_left_out[0:95]),
		.chanx_right_out(cbx_2__1__4_chanx_right_out[0:95]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_f2a_i_0_(cbx_2__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_f2a_i_0_(cbx_2__1__4_bottom_grid_top_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_f2a_i_0_(cbx_2__1__4_bottom_grid_top_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_f2a_i_0_(cbx_2__1__4_bottom_grid_top_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_f2a_i_0_(cbx_2__1__4_bottom_grid_top_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_f2a_i_0_(cbx_2__1__4_bottom_grid_top_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_f2a_i_0_(cbx_2__1__4_bottom_grid_top_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_f2a_i_0_(cbx_2__1__4_bottom_grid_top_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_f2a_i_0_(cbx_2__1__4_bottom_grid_top_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_9__pin_f2a_i_0_(cbx_2__1__4_bottom_grid_top_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_10__pin_f2a_i_0_(cbx_2__1__4_bottom_grid_top_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_11__pin_f2a_i_0_(cbx_2__1__4_bottom_grid_top_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_12__pin_f2a_i_0_(cbx_2__1__4_bottom_grid_top_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_13__pin_f2a_i_0_(cbx_2__1__4_bottom_grid_top_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_14__pin_f2a_i_0_(cbx_2__1__4_bottom_grid_top_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_15__pin_f2a_i_0_(cbx_2__1__4_bottom_grid_top_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_16__pin_f2a_i_0_(cbx_2__1__4_bottom_grid_top_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_17__pin_f2a_i_0_(cbx_2__1__4_bottom_grid_top_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_18__pin_f2a_i_0_(cbx_2__1__4_bottom_grid_top_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_19__pin_f2a_i_0_(cbx_2__1__4_bottom_grid_top_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.ccff_tail(cbx_2__1__4_ccff_tail));

	cbx_2__1_ cbx_9__1_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chanx_left_in(sb_2__1__3_chanx_right_out[0:95]),
		.chanx_right_in(sb_9__1__0_chanx_left_out[0:95]),
		.ccff_head(sb_9__1__0_ccff_tail),
		.chanx_left_out(cbx_2__1__5_chanx_left_out[0:95]),
		.chanx_right_out(cbx_2__1__5_chanx_right_out[0:95]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_f2a_i_0_(cbx_2__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_f2a_i_0_(cbx_2__1__5_bottom_grid_top_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_f2a_i_0_(cbx_2__1__5_bottom_grid_top_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_f2a_i_0_(cbx_2__1__5_bottom_grid_top_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_f2a_i_0_(cbx_2__1__5_bottom_grid_top_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_f2a_i_0_(cbx_2__1__5_bottom_grid_top_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_f2a_i_0_(cbx_2__1__5_bottom_grid_top_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_f2a_i_0_(cbx_2__1__5_bottom_grid_top_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_f2a_i_0_(cbx_2__1__5_bottom_grid_top_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_9__pin_f2a_i_0_(cbx_2__1__5_bottom_grid_top_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_10__pin_f2a_i_0_(cbx_2__1__5_bottom_grid_top_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_11__pin_f2a_i_0_(cbx_2__1__5_bottom_grid_top_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_12__pin_f2a_i_0_(cbx_2__1__5_bottom_grid_top_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_13__pin_f2a_i_0_(cbx_2__1__5_bottom_grid_top_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_14__pin_f2a_i_0_(cbx_2__1__5_bottom_grid_top_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_15__pin_f2a_i_0_(cbx_2__1__5_bottom_grid_top_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_16__pin_f2a_i_0_(cbx_2__1__5_bottom_grid_top_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_17__pin_f2a_i_0_(cbx_2__1__5_bottom_grid_top_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_18__pin_f2a_i_0_(cbx_2__1__5_bottom_grid_top_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_19__pin_f2a_i_0_(cbx_2__1__5_bottom_grid_top_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.ccff_tail(cbx_2__1__5_ccff_tail));

	cbx_2__2_ cbx_2__2_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chanx_left_in(sb_1__2__0_chanx_right_out[0:95]),
		.chanx_right_in(sb_2__2__0_chanx_left_out[0:95]),
		.ccff_head(sb_2__2__0_ccff_tail),
		.chanx_left_out(cbx_2__2__0_chanx_left_out[0:95]),
		.chanx_right_out(cbx_2__2__0_chanx_right_out[0:95]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.ccff_tail(cbx_2__2__0_ccff_tail));

	cbx_2__2_ cbx_2__3_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chanx_left_in(sb_1__2__1_chanx_right_out[0:95]),
		.chanx_right_in(sb_2__2__1_chanx_left_out[0:95]),
		.ccff_head(sb_2__2__1_ccff_tail),
		.chanx_left_out(cbx_2__2__1_chanx_left_out[0:95]),
		.chanx_right_out(cbx_2__2__1_chanx_right_out[0:95]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.ccff_tail(ccff_tail[4]));

	cbx_2__2_ cbx_2__4_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chanx_left_in(sb_1__2__2_chanx_right_out[0:95]),
		.chanx_right_in(sb_2__2__2_chanx_left_out[0:95]),
		.ccff_head(sb_2__2__2_ccff_tail),
		.chanx_left_out(cbx_2__2__2_chanx_left_out[0:95]),
		.chanx_right_out(cbx_2__2__2_chanx_right_out[0:95]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.ccff_tail(cbx_2__2__2_ccff_tail));

	cbx_2__2_ cbx_2__5_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chanx_left_in(sb_1__2__3_chanx_right_out[0:95]),
		.chanx_right_in(sb_2__2__3_chanx_left_out[0:95]),
		.ccff_head(sb_2__2__3_ccff_tail),
		.chanx_left_out(cbx_2__2__3_chanx_left_out[0:95]),
		.chanx_right_out(cbx_2__2__3_chanx_right_out[0:95]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.ccff_tail(cbx_2__2__3_ccff_tail));

	cbx_2__2_ cbx_2__6_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chanx_left_in(sb_1__2__4_chanx_right_out[0:95]),
		.chanx_right_in(sb_2__2__4_chanx_left_out[0:95]),
		.ccff_head(sb_2__2__4_ccff_tail),
		.chanx_left_out(cbx_2__2__4_chanx_left_out[0:95]),
		.chanx_right_out(cbx_2__2__4_chanx_right_out[0:95]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.ccff_tail(cbx_2__2__4_ccff_tail));

	cbx_2__2_ cbx_3__2_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chanx_left_in(sb_2__2__0_chanx_right_out[0:95]),
		.chanx_right_in(sb_3__2__0_chanx_left_out[0:95]),
		.ccff_head(sb_3__2__0_ccff_tail),
		.chanx_left_out(cbx_2__2__5_chanx_left_out[0:95]),
		.chanx_right_out(cbx_2__2__5_chanx_right_out[0:95]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.ccff_tail(cbx_2__2__5_ccff_tail));

	cbx_2__2_ cbx_3__3_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chanx_left_in(sb_2__2__1_chanx_right_out[0:95]),
		.chanx_right_in(sb_3__2__1_chanx_left_out[0:95]),
		.ccff_head(sb_3__2__1_ccff_tail),
		.chanx_left_out(cbx_2__2__6_chanx_left_out[0:95]),
		.chanx_right_out(cbx_2__2__6_chanx_right_out[0:95]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__6_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.ccff_tail(cbx_2__2__6_ccff_tail));

	cbx_2__2_ cbx_3__4_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chanx_left_in(sb_2__2__2_chanx_right_out[0:95]),
		.chanx_right_in(sb_3__4__0_chanx_left_out[0:95]),
		.ccff_head(sb_3__4__0_ccff_tail),
		.chanx_left_out(cbx_2__2__7_chanx_left_out[0:95]),
		.chanx_right_out(cbx_2__2__7_chanx_right_out[0:95]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__7_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.ccff_tail(cbx_2__2__7_ccff_tail));

	cbx_2__2_ cbx_3__5_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chanx_left_in(sb_2__2__3_chanx_right_out[0:95]),
		.chanx_right_in(sb_3__2__2_chanx_left_out[0:95]),
		.ccff_head(sb_3__2__2_ccff_tail),
		.chanx_left_out(cbx_2__2__8_chanx_left_out[0:95]),
		.chanx_right_out(cbx_2__2__8_chanx_right_out[0:95]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__8_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.ccff_tail(cbx_2__2__8_ccff_tail));

	cbx_2__2_ cbx_3__6_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chanx_left_in(sb_2__2__4_chanx_right_out[0:95]),
		.chanx_right_in(sb_3__2__3_chanx_left_out[0:95]),
		.ccff_head(ccff_head[8]),
		.chanx_left_out(cbx_2__2__9_chanx_left_out[0:95]),
		.chanx_right_out(cbx_2__2__9_chanx_right_out[0:95]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__9_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.ccff_tail(cbx_2__2__9_ccff_tail));

	cbx_2__2_ cbx_5__2_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chanx_left_in(sb_4__2__0_chanx_right_out[0:95]),
		.chanx_right_in(sb_2__2__5_chanx_left_out[0:95]),
		.ccff_head(sb_2__2__5_ccff_tail),
		.chanx_left_out(cbx_2__2__10_chanx_left_out[0:95]),
		.chanx_right_out(cbx_2__2__10_chanx_right_out[0:95]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__10_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.ccff_tail(cbx_2__2__10_ccff_tail));

	cbx_2__2_ cbx_5__3_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chanx_left_in(sb_4__3__0_chanx_right_out[0:95]),
		.chanx_right_in(sb_2__2__6_chanx_left_out[0:95]),
		.ccff_head(sb_2__2__6_ccff_tail),
		.chanx_left_out(cbx_2__2__11_chanx_left_out[0:95]),
		.chanx_right_out(cbx_2__2__11_chanx_right_out[0:95]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__11_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.ccff_tail(cbx_2__2__11_ccff_tail));

	cbx_2__2_ cbx_5__4_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chanx_left_in(sb_4__4__0_chanx_right_out[0:95]),
		.chanx_right_in(sb_2__2__7_chanx_left_out[0:95]),
		.ccff_head(sb_2__2__7_ccff_tail),
		.chanx_left_out(cbx_2__2__12_chanx_left_out[0:95]),
		.chanx_right_out(cbx_2__2__12_chanx_right_out[0:95]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__12_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.ccff_tail(cbx_2__2__12_ccff_tail));

	cbx_2__2_ cbx_5__5_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chanx_left_in(sb_4__2__1_chanx_right_out[0:95]),
		.chanx_right_in(sb_2__2__8_chanx_left_out[0:95]),
		.ccff_head(sb_2__2__8_ccff_tail),
		.chanx_left_out(cbx_2__2__13_chanx_left_out[0:95]),
		.chanx_right_out(cbx_2__2__13_chanx_right_out[0:95]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__13_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.ccff_tail(cbx_2__2__13_ccff_tail));

	cbx_2__2_ cbx_5__6_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chanx_left_in(sb_4__3__1_chanx_right_out[0:95]),
		.chanx_right_in(sb_2__2__9_chanx_left_out[0:95]),
		.ccff_head(sb_2__2__9_ccff_tail),
		.chanx_left_out(cbx_2__2__14_chanx_left_out[0:95]),
		.chanx_right_out(cbx_2__2__14_chanx_right_out[0:95]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__14_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.ccff_tail(cbx_2__2__14_ccff_tail));

	cbx_2__2_ cbx_6__2_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chanx_left_in(sb_2__2__5_chanx_right_out[0:95]),
		.chanx_right_in(sb_3__2__4_chanx_left_out[0:95]),
		.ccff_head(sb_3__2__4_ccff_tail),
		.chanx_left_out(cbx_2__2__15_chanx_left_out[0:95]),
		.chanx_right_out(cbx_2__2__15_chanx_right_out[0:95]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__15_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.ccff_tail(cbx_2__2__15_ccff_tail));

	cbx_2__2_ cbx_6__3_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chanx_left_in(sb_2__2__6_chanx_right_out[0:95]),
		.chanx_right_in(sb_3__2__5_chanx_left_out[0:95]),
		.ccff_head(sb_3__2__5_ccff_tail),
		.chanx_left_out(cbx_2__2__16_chanx_left_out[0:95]),
		.chanx_right_out(cbx_2__2__16_chanx_right_out[0:95]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__16_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.ccff_tail(cbx_2__2__16_ccff_tail));

	cbx_2__2_ cbx_6__4_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chanx_left_in(sb_2__2__7_chanx_right_out[0:95]),
		.chanx_right_in(sb_3__2__6_chanx_left_out[0:95]),
		.ccff_head(sb_3__2__6_ccff_tail),
		.chanx_left_out(cbx_2__2__17_chanx_left_out[0:95]),
		.chanx_right_out(cbx_2__2__17_chanx_right_out[0:95]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__17_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.ccff_tail(cbx_2__2__17_ccff_tail));

	cbx_2__2_ cbx_6__5_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chanx_left_in(sb_2__2__8_chanx_right_out[0:95]),
		.chanx_right_in(sb_3__2__7_chanx_left_out[0:95]),
		.ccff_head(sb_3__2__7_ccff_tail),
		.chanx_left_out(cbx_2__2__18_chanx_left_out[0:95]),
		.chanx_right_out(cbx_2__2__18_chanx_right_out[0:95]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__18_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.ccff_tail(ccff_tail[6]));

	cbx_2__2_ cbx_6__6_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chanx_left_in(sb_2__2__9_chanx_right_out[0:95]),
		.chanx_right_in(sb_3__2__8_chanx_left_out[0:95]),
		.ccff_head(sb_3__2__8_ccff_tail),
		.chanx_left_out(cbx_2__2__19_chanx_left_out[0:95]),
		.chanx_right_out(cbx_2__2__19_chanx_right_out[0:95]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__19_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.ccff_tail(cbx_2__2__19_ccff_tail));

	cbx_2__2_ cbx_8__2_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chanx_left_in(sb_7__2__0_chanx_right_out[0:95]),
		.chanx_right_in(sb_2__2__10_chanx_left_out[0:95]),
		.ccff_head(sb_2__2__10_ccff_tail),
		.chanx_left_out(cbx_2__2__20_chanx_left_out[0:95]),
		.chanx_right_out(cbx_2__2__20_chanx_right_out[0:95]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__20_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.ccff_tail(cbx_2__2__20_ccff_tail));

	cbx_2__2_ cbx_8__3_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chanx_left_in(sb_7__2__1_chanx_right_out[0:95]),
		.chanx_right_in(sb_2__2__11_chanx_left_out[0:95]),
		.ccff_head(sb_2__2__11_ccff_tail),
		.chanx_left_out(cbx_2__2__21_chanx_left_out[0:95]),
		.chanx_right_out(cbx_2__2__21_chanx_right_out[0:95]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__21_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.ccff_tail(cbx_2__2__21_ccff_tail));

	cbx_2__2_ cbx_8__4_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chanx_left_in(sb_7__2__2_chanx_right_out[0:95]),
		.chanx_right_in(sb_2__2__12_chanx_left_out[0:95]),
		.ccff_head(sb_2__2__12_ccff_tail),
		.chanx_left_out(cbx_2__2__22_chanx_left_out[0:95]),
		.chanx_right_out(cbx_2__2__22_chanx_right_out[0:95]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__22_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.ccff_tail(cbx_2__2__22_ccff_tail));

	cbx_2__2_ cbx_8__5_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chanx_left_in(sb_7__2__3_chanx_right_out[0:95]),
		.chanx_right_in(sb_2__2__13_chanx_left_out[0:95]),
		.ccff_head(sb_2__2__13_ccff_tail),
		.chanx_left_out(cbx_2__2__23_chanx_left_out[0:95]),
		.chanx_right_out(cbx_2__2__23_chanx_right_out[0:95]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__23_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.ccff_tail(cbx_2__2__23_ccff_tail));

	cbx_2__2_ cbx_8__6_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chanx_left_in(sb_7__2__4_chanx_right_out[0:95]),
		.chanx_right_in(sb_2__2__14_chanx_left_out[0:95]),
		.ccff_head(sb_2__2__14_ccff_tail),
		.chanx_left_out(cbx_2__2__24_chanx_left_out[0:95]),
		.chanx_right_out(cbx_2__2__24_chanx_right_out[0:95]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__24_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.ccff_tail(cbx_2__2__24_ccff_tail));

	cbx_2__2_ cbx_9__2_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chanx_left_in(sb_2__2__10_chanx_right_out[0:95]),
		.chanx_right_in(sb_9__2__0_chanx_left_out[0:95]),
		.ccff_head(sb_9__2__0_ccff_tail),
		.chanx_left_out(cbx_2__2__25_chanx_left_out[0:95]),
		.chanx_right_out(cbx_2__2__25_chanx_right_out[0:95]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__25_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.ccff_tail(cbx_2__2__25_ccff_tail));

	cbx_2__2_ cbx_9__3_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chanx_left_in(sb_2__2__11_chanx_right_out[0:95]),
		.chanx_right_in(sb_9__2__1_chanx_left_out[0:95]),
		.ccff_head(sb_9__2__1_ccff_tail),
		.chanx_left_out(cbx_2__2__26_chanx_left_out[0:95]),
		.chanx_right_out(cbx_2__2__26_chanx_right_out[0:95]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__26_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.ccff_tail(cbx_2__2__26_ccff_tail));

	cbx_2__2_ cbx_9__4_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chanx_left_in(sb_2__2__12_chanx_right_out[0:95]),
		.chanx_right_in(sb_9__2__2_chanx_left_out[0:95]),
		.ccff_head(sb_9__2__2_ccff_tail),
		.chanx_left_out(cbx_2__2__27_chanx_left_out[0:95]),
		.chanx_right_out(cbx_2__2__27_chanx_right_out[0:95]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__27_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.ccff_tail(cbx_2__2__27_ccff_tail));

	cbx_2__2_ cbx_9__5_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chanx_left_in(sb_2__2__13_chanx_right_out[0:95]),
		.chanx_right_in(sb_9__2__3_chanx_left_out[0:95]),
		.ccff_head(sb_9__2__3_ccff_tail),
		.chanx_left_out(cbx_2__2__28_chanx_left_out[0:95]),
		.chanx_right_out(cbx_2__2__28_chanx_right_out[0:95]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__28_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.ccff_tail(cbx_2__2__28_ccff_tail));

	cbx_2__2_ cbx_9__6_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chanx_left_in(sb_2__2__14_chanx_right_out[0:95]),
		.chanx_right_in(sb_9__2__4_chanx_left_out[0:95]),
		.ccff_head(sb_9__2__4_ccff_tail),
		.chanx_left_out(cbx_2__2__29_chanx_left_out[0:95]),
		.chanx_right_out(cbx_2__2__29_chanx_right_out[0:95]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__2__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__2__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__2__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__2__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__2__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__2__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__2__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__2__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__2__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__2__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__2__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__2__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__2__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__2__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__2__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__2__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__2__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__2__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__2__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__2__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__2__29_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.ccff_tail(cbx_2__2__29_ccff_tail));

	cbx_2__7_ cbx_2__7_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chanx_left_in(sb_1__7__0_chanx_right_out[0:95]),
		.chanx_right_in(sb_2__7__0_chanx_left_out[0:95]),
		.ccff_head(sb_2__7__0_ccff_tail),
		.chanx_left_out(cbx_2__7__0_chanx_left_out[0:95]),
		.chanx_right_out(cbx_2__7__0_chanx_right_out[0:95]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_f2a_i_0_(cbx_2__7__0_top_grid_bottom_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_f2a_i_0_(cbx_2__7__0_top_grid_bottom_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_f2a_i_0_(cbx_2__7__0_top_grid_bottom_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_f2a_i_0_(cbx_2__7__0_top_grid_bottom_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_f2a_i_0_(cbx_2__7__0_top_grid_bottom_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_f2a_i_0_(cbx_2__7__0_top_grid_bottom_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_f2a_i_0_(cbx_2__7__0_top_grid_bottom_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_f2a_i_0_(cbx_2__7__0_top_grid_bottom_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_8__pin_f2a_i_0_(cbx_2__7__0_top_grid_bottom_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_9__pin_f2a_i_0_(cbx_2__7__0_top_grid_bottom_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_10__pin_f2a_i_0_(cbx_2__7__0_top_grid_bottom_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_11__pin_f2a_i_0_(cbx_2__7__0_top_grid_bottom_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_12__pin_f2a_i_0_(cbx_2__7__0_top_grid_bottom_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_13__pin_f2a_i_0_(cbx_2__7__0_top_grid_bottom_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_14__pin_f2a_i_0_(cbx_2__7__0_top_grid_bottom_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_15__pin_f2a_i_0_(cbx_2__7__0_top_grid_bottom_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_16__pin_f2a_i_0_(cbx_2__7__0_top_grid_bottom_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_17__pin_f2a_i_0_(cbx_2__7__0_top_grid_bottom_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_18__pin_f2a_i_0_(cbx_2__7__0_top_grid_bottom_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_19__pin_f2a_i_0_(cbx_2__7__0_top_grid_bottom_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__7__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__7__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__7__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__7__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__7__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__7__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__7__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__7__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__7__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__7__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__7__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__7__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__7__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__7__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__7__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__7__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__7__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__7__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__7__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__7__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__7__0_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.ccff_tail(cbx_2__7__0_ccff_tail));

	cbx_2__7_ cbx_3__7_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chanx_left_in(sb_2__7__0_chanx_right_out[0:95]),
		.chanx_right_in(sb_3__7__0_chanx_left_out[0:95]),
		.ccff_head(sb_3__7__0_ccff_tail),
		.chanx_left_out(cbx_2__7__1_chanx_left_out[0:95]),
		.chanx_right_out(cbx_2__7__1_chanx_right_out[0:95]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_f2a_i_0_(cbx_2__7__1_top_grid_bottom_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_f2a_i_0_(cbx_2__7__1_top_grid_bottom_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_f2a_i_0_(cbx_2__7__1_top_grid_bottom_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_f2a_i_0_(cbx_2__7__1_top_grid_bottom_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_f2a_i_0_(cbx_2__7__1_top_grid_bottom_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_f2a_i_0_(cbx_2__7__1_top_grid_bottom_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_f2a_i_0_(cbx_2__7__1_top_grid_bottom_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_f2a_i_0_(cbx_2__7__1_top_grid_bottom_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_8__pin_f2a_i_0_(cbx_2__7__1_top_grid_bottom_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_9__pin_f2a_i_0_(cbx_2__7__1_top_grid_bottom_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_10__pin_f2a_i_0_(cbx_2__7__1_top_grid_bottom_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_11__pin_f2a_i_0_(cbx_2__7__1_top_grid_bottom_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_12__pin_f2a_i_0_(cbx_2__7__1_top_grid_bottom_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_13__pin_f2a_i_0_(cbx_2__7__1_top_grid_bottom_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_14__pin_f2a_i_0_(cbx_2__7__1_top_grid_bottom_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_15__pin_f2a_i_0_(cbx_2__7__1_top_grid_bottom_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_16__pin_f2a_i_0_(cbx_2__7__1_top_grid_bottom_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_17__pin_f2a_i_0_(cbx_2__7__1_top_grid_bottom_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_18__pin_f2a_i_0_(cbx_2__7__1_top_grid_bottom_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_19__pin_f2a_i_0_(cbx_2__7__1_top_grid_bottom_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__7__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__7__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__7__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__7__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__7__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__7__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__7__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__7__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__7__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__7__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__7__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__7__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__7__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__7__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__7__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__7__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__7__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__7__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__7__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__7__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__7__1_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.ccff_tail(cbx_2__7__1_ccff_tail));

	cbx_2__7_ cbx_5__7_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chanx_left_in(sb_4__7__0_chanx_right_out[0:95]),
		.chanx_right_in(sb_2__7__1_chanx_left_out[0:95]),
		.ccff_head(sb_2__7__1_ccff_tail),
		.chanx_left_out(cbx_2__7__2_chanx_left_out[0:95]),
		.chanx_right_out(cbx_2__7__2_chanx_right_out[0:95]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_f2a_i_0_(cbx_2__7__2_top_grid_bottom_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_f2a_i_0_(cbx_2__7__2_top_grid_bottom_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_f2a_i_0_(cbx_2__7__2_top_grid_bottom_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_f2a_i_0_(cbx_2__7__2_top_grid_bottom_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_f2a_i_0_(cbx_2__7__2_top_grid_bottom_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_f2a_i_0_(cbx_2__7__2_top_grid_bottom_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_f2a_i_0_(cbx_2__7__2_top_grid_bottom_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_f2a_i_0_(cbx_2__7__2_top_grid_bottom_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_8__pin_f2a_i_0_(cbx_2__7__2_top_grid_bottom_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_9__pin_f2a_i_0_(cbx_2__7__2_top_grid_bottom_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_10__pin_f2a_i_0_(cbx_2__7__2_top_grid_bottom_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_11__pin_f2a_i_0_(cbx_2__7__2_top_grid_bottom_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_12__pin_f2a_i_0_(cbx_2__7__2_top_grid_bottom_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_13__pin_f2a_i_0_(cbx_2__7__2_top_grid_bottom_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_14__pin_f2a_i_0_(cbx_2__7__2_top_grid_bottom_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_15__pin_f2a_i_0_(cbx_2__7__2_top_grid_bottom_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_16__pin_f2a_i_0_(cbx_2__7__2_top_grid_bottom_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_17__pin_f2a_i_0_(cbx_2__7__2_top_grid_bottom_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_18__pin_f2a_i_0_(cbx_2__7__2_top_grid_bottom_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_19__pin_f2a_i_0_(cbx_2__7__2_top_grid_bottom_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__7__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__7__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__7__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__7__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__7__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__7__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__7__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__7__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__7__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__7__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__7__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__7__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__7__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__7__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__7__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__7__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__7__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__7__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__7__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__7__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__7__2_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.ccff_tail(cbx_2__7__2_ccff_tail));

	cbx_2__7_ cbx_6__7_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chanx_left_in(sb_2__7__1_chanx_right_out[0:95]),
		.chanx_right_in(sb_3__7__1_chanx_left_out[0:95]),
		.ccff_head(sb_3__7__1_ccff_tail),
		.chanx_left_out(cbx_2__7__3_chanx_left_out[0:95]),
		.chanx_right_out(cbx_2__7__3_chanx_right_out[0:95]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_f2a_i_0_(cbx_2__7__3_top_grid_bottom_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_f2a_i_0_(cbx_2__7__3_top_grid_bottom_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_f2a_i_0_(cbx_2__7__3_top_grid_bottom_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_f2a_i_0_(cbx_2__7__3_top_grid_bottom_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_f2a_i_0_(cbx_2__7__3_top_grid_bottom_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_f2a_i_0_(cbx_2__7__3_top_grid_bottom_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_f2a_i_0_(cbx_2__7__3_top_grid_bottom_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_f2a_i_0_(cbx_2__7__3_top_grid_bottom_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_8__pin_f2a_i_0_(cbx_2__7__3_top_grid_bottom_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_9__pin_f2a_i_0_(cbx_2__7__3_top_grid_bottom_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_10__pin_f2a_i_0_(cbx_2__7__3_top_grid_bottom_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_11__pin_f2a_i_0_(cbx_2__7__3_top_grid_bottom_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_12__pin_f2a_i_0_(cbx_2__7__3_top_grid_bottom_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_13__pin_f2a_i_0_(cbx_2__7__3_top_grid_bottom_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_14__pin_f2a_i_0_(cbx_2__7__3_top_grid_bottom_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_15__pin_f2a_i_0_(cbx_2__7__3_top_grid_bottom_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_16__pin_f2a_i_0_(cbx_2__7__3_top_grid_bottom_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_17__pin_f2a_i_0_(cbx_2__7__3_top_grid_bottom_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_18__pin_f2a_i_0_(cbx_2__7__3_top_grid_bottom_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_19__pin_f2a_i_0_(cbx_2__7__3_top_grid_bottom_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__7__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__7__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__7__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__7__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__7__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__7__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__7__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__7__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__7__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__7__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__7__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__7__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__7__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__7__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__7__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__7__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__7__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__7__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__7__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__7__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__7__3_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.ccff_tail(cbx_2__7__3_ccff_tail));

	cbx_2__7_ cbx_8__7_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chanx_left_in(sb_7__7__0_chanx_right_out[0:95]),
		.chanx_right_in(sb_2__7__2_chanx_left_out[0:95]),
		.ccff_head(sb_2__7__2_ccff_tail),
		.chanx_left_out(cbx_2__7__4_chanx_left_out[0:95]),
		.chanx_right_out(cbx_2__7__4_chanx_right_out[0:95]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_f2a_i_0_(cbx_2__7__4_top_grid_bottom_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_f2a_i_0_(cbx_2__7__4_top_grid_bottom_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_f2a_i_0_(cbx_2__7__4_top_grid_bottom_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_f2a_i_0_(cbx_2__7__4_top_grid_bottom_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_f2a_i_0_(cbx_2__7__4_top_grid_bottom_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_f2a_i_0_(cbx_2__7__4_top_grid_bottom_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_f2a_i_0_(cbx_2__7__4_top_grid_bottom_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_f2a_i_0_(cbx_2__7__4_top_grid_bottom_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_8__pin_f2a_i_0_(cbx_2__7__4_top_grid_bottom_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_9__pin_f2a_i_0_(cbx_2__7__4_top_grid_bottom_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_10__pin_f2a_i_0_(cbx_2__7__4_top_grid_bottom_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_11__pin_f2a_i_0_(cbx_2__7__4_top_grid_bottom_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_12__pin_f2a_i_0_(cbx_2__7__4_top_grid_bottom_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_13__pin_f2a_i_0_(cbx_2__7__4_top_grid_bottom_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_14__pin_f2a_i_0_(cbx_2__7__4_top_grid_bottom_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_15__pin_f2a_i_0_(cbx_2__7__4_top_grid_bottom_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_16__pin_f2a_i_0_(cbx_2__7__4_top_grid_bottom_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_17__pin_f2a_i_0_(cbx_2__7__4_top_grid_bottom_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_18__pin_f2a_i_0_(cbx_2__7__4_top_grid_bottom_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_19__pin_f2a_i_0_(cbx_2__7__4_top_grid_bottom_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__7__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__7__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__7__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__7__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__7__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__7__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__7__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__7__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__7__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__7__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__7__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__7__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__7__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__7__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__7__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__7__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__7__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__7__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__7__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__7__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__7__4_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.ccff_tail(cbx_2__7__4_ccff_tail));

	cbx_2__7_ cbx_9__7_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chanx_left_in(sb_2__7__2_chanx_right_out[0:95]),
		.chanx_right_in(sb_9__7__0_chanx_left_out[0:95]),
		.ccff_head(sb_9__7__0_ccff_tail),
		.chanx_left_out(cbx_2__7__5_chanx_left_out[0:95]),
		.chanx_right_out(cbx_2__7__5_chanx_right_out[0:95]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_f2a_i_0_(cbx_2__7__5_top_grid_bottom_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_f2a_i_0_(cbx_2__7__5_top_grid_bottom_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_f2a_i_0_(cbx_2__7__5_top_grid_bottom_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_f2a_i_0_(cbx_2__7__5_top_grid_bottom_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_f2a_i_0_(cbx_2__7__5_top_grid_bottom_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_f2a_i_0_(cbx_2__7__5_top_grid_bottom_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_f2a_i_0_(cbx_2__7__5_top_grid_bottom_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_f2a_i_0_(cbx_2__7__5_top_grid_bottom_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_8__pin_f2a_i_0_(cbx_2__7__5_top_grid_bottom_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_9__pin_f2a_i_0_(cbx_2__7__5_top_grid_bottom_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_10__pin_f2a_i_0_(cbx_2__7__5_top_grid_bottom_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_11__pin_f2a_i_0_(cbx_2__7__5_top_grid_bottom_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_12__pin_f2a_i_0_(cbx_2__7__5_top_grid_bottom_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_13__pin_f2a_i_0_(cbx_2__7__5_top_grid_bottom_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_14__pin_f2a_i_0_(cbx_2__7__5_top_grid_bottom_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_15__pin_f2a_i_0_(cbx_2__7__5_top_grid_bottom_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_16__pin_f2a_i_0_(cbx_2__7__5_top_grid_bottom_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_17__pin_f2a_i_0_(cbx_2__7__5_top_grid_bottom_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_18__pin_f2a_i_0_(cbx_2__7__5_top_grid_bottom_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_19__pin_f2a_i_0_(cbx_2__7__5_top_grid_bottom_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_2__7__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_2__7__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_(cbx_2__7__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_(cbx_2__7__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_(cbx_2__7__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_(cbx_2__7__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_(cbx_2__7__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_(cbx_2__7__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_(cbx_2__7__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_(cbx_2__7__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_2__7__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_2__7__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_(cbx_2__7__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_(cbx_2__7__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_(cbx_2__7__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_(cbx_2__7__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_(cbx_2__7__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_(cbx_2__7__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_(cbx_2__7__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_(cbx_2__7__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_(cbx_2__7__5_bottom_grid_top_width_0_height_0_subtile_0__pin_cin_trick_0_),
		.ccff_tail(cbx_2__7__5_ccff_tail));

	cbx_4__1_ cbx_4__1_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chanx_left_in(sb_3__1__0_chanx_right_out[0:95]),
		.chanx_right_in(sb_4__1__0_chanx_left_out[0:95]),
		.ccff_head(sb_4__1__0_ccff_tail),
		.chanx_left_out(cbx_4__1__0_chanx_left_out[0:95]),
		.chanx_right_out(cbx_4__1__0_chanx_right_out[0:95]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_a_i_0_(cbx_4__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_a_i_1_(cbx_4__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_a_i_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_acc_fir_i_0_(cbx_4__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_acc_fir_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_lreset_0_(cbx_4__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_lreset_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_feedback_0_(cbx_4__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_feedback_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_feedback_1_(cbx_4__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_feedback_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_feedback_2_(cbx_4__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_feedback_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_shift_right_0_(cbx_4__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_shift_right_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_shift_right_1_(cbx_4__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_shift_right_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_shift_right_2_(cbx_4__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_shift_right_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_shift_right_3_(cbx_4__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_shift_right_3_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_shift_right_4_(cbx_4__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_shift_right_4_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_shift_right_5_(cbx_4__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_shift_right_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_f2a_i_0_(cbx_4__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_f2a_i_0_(cbx_4__1__0_bottom_grid_top_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_f2a_i_0_(cbx_4__1__0_bottom_grid_top_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_f2a_i_0_(cbx_4__1__0_bottom_grid_top_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_f2a_i_0_(cbx_4__1__0_bottom_grid_top_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_f2a_i_0_(cbx_4__1__0_bottom_grid_top_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_f2a_i_0_(cbx_4__1__0_bottom_grid_top_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_f2a_i_0_(cbx_4__1__0_bottom_grid_top_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_f2a_i_0_(cbx_4__1__0_bottom_grid_top_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_9__pin_f2a_i_0_(cbx_4__1__0_bottom_grid_top_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_10__pin_f2a_i_0_(cbx_4__1__0_bottom_grid_top_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_11__pin_f2a_i_0_(cbx_4__1__0_bottom_grid_top_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_12__pin_f2a_i_0_(cbx_4__1__0_bottom_grid_top_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_13__pin_f2a_i_0_(cbx_4__1__0_bottom_grid_top_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_14__pin_f2a_i_0_(cbx_4__1__0_bottom_grid_top_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_15__pin_f2a_i_0_(cbx_4__1__0_bottom_grid_top_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_16__pin_f2a_i_0_(cbx_4__1__0_bottom_grid_top_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_17__pin_f2a_i_0_(cbx_4__1__0_bottom_grid_top_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_18__pin_f2a_i_0_(cbx_4__1__0_bottom_grid_top_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_19__pin_f2a_i_0_(cbx_4__1__0_bottom_grid_top_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.ccff_tail(cbx_4__1__0_ccff_tail));

	cbx_4__4_ cbx_4__4_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chanx_left_in(sb_3__4__0_chanx_right_out[0:95]),
		.chanx_right_in(sb_4__4__0_chanx_left_out[0:95]),
		.ccff_head(sb_4__4__0_ccff_tail),
		.chanx_left_out(cbx_4__4__0_chanx_left_out[0:95]),
		.chanx_right_out(cbx_4__4__0_chanx_right_out[0:95]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_a_i_0_(cbx_4__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_a_i_1_(cbx_4__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_a_i_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_acc_fir_i_0_(cbx_4__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_acc_fir_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_lreset_0_(cbx_4__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_lreset_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_feedback_0_(cbx_4__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_feedback_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_feedback_1_(cbx_4__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_feedback_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_feedback_2_(cbx_4__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_feedback_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_shift_right_0_(cbx_4__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_shift_right_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_shift_right_1_(cbx_4__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_shift_right_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_shift_right_2_(cbx_4__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_shift_right_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_shift_right_3_(cbx_4__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_shift_right_3_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_shift_right_4_(cbx_4__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_shift_right_4_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_shift_right_5_(cbx_4__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_shift_right_5_),
		.ccff_tail(cbx_4__4__0_ccff_tail));

	cbx_4__7_ cbx_4__7_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chanx_left_in(sb_3__7__0_chanx_right_out[0:95]),
		.chanx_right_in(sb_4__7__0_chanx_left_out[0:95]),
		.ccff_head(sb_4__7__0_ccff_tail),
		.chanx_left_out(cbx_4__7__0_chanx_left_out[0:95]),
		.chanx_right_out(cbx_4__7__0_chanx_right_out[0:95]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_f2a_i_0_(cbx_4__7__0_top_grid_bottom_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_f2a_i_0_(cbx_4__7__0_top_grid_bottom_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_f2a_i_0_(cbx_4__7__0_top_grid_bottom_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_f2a_i_0_(cbx_4__7__0_top_grid_bottom_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_f2a_i_0_(cbx_4__7__0_top_grid_bottom_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_f2a_i_0_(cbx_4__7__0_top_grid_bottom_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_f2a_i_0_(cbx_4__7__0_top_grid_bottom_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_f2a_i_0_(cbx_4__7__0_top_grid_bottom_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_8__pin_f2a_i_0_(cbx_4__7__0_top_grid_bottom_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_9__pin_f2a_i_0_(cbx_4__7__0_top_grid_bottom_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_10__pin_f2a_i_0_(cbx_4__7__0_top_grid_bottom_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_11__pin_f2a_i_0_(cbx_4__7__0_top_grid_bottom_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_12__pin_f2a_i_0_(cbx_4__7__0_top_grid_bottom_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_13__pin_f2a_i_0_(cbx_4__7__0_top_grid_bottom_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_14__pin_f2a_i_0_(cbx_4__7__0_top_grid_bottom_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_15__pin_f2a_i_0_(cbx_4__7__0_top_grid_bottom_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_16__pin_f2a_i_0_(cbx_4__7__0_top_grid_bottom_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_17__pin_f2a_i_0_(cbx_4__7__0_top_grid_bottom_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_18__pin_f2a_i_0_(cbx_4__7__0_top_grid_bottom_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_19__pin_f2a_i_0_(cbx_4__7__0_top_grid_bottom_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.ccff_tail(cbx_4__7__0_ccff_tail));

	cbx_4__7_ cbx_7__7_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chanx_left_in(sb_3__7__1_chanx_right_out[0:95]),
		.chanx_right_in(sb_7__7__0_chanx_left_out[0:95]),
		.ccff_head(sb_7__7__0_ccff_tail),
		.chanx_left_out(cbx_4__7__1_chanx_left_out[0:95]),
		.chanx_right_out(cbx_4__7__1_chanx_right_out[0:95]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_f2a_i_0_(cbx_4__7__1_top_grid_bottom_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_f2a_i_0_(cbx_4__7__1_top_grid_bottom_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_f2a_i_0_(cbx_4__7__1_top_grid_bottom_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_f2a_i_0_(cbx_4__7__1_top_grid_bottom_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_f2a_i_0_(cbx_4__7__1_top_grid_bottom_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_f2a_i_0_(cbx_4__7__1_top_grid_bottom_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_f2a_i_0_(cbx_4__7__1_top_grid_bottom_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_f2a_i_0_(cbx_4__7__1_top_grid_bottom_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_8__pin_f2a_i_0_(cbx_4__7__1_top_grid_bottom_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_9__pin_f2a_i_0_(cbx_4__7__1_top_grid_bottom_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_10__pin_f2a_i_0_(cbx_4__7__1_top_grid_bottom_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_11__pin_f2a_i_0_(cbx_4__7__1_top_grid_bottom_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_12__pin_f2a_i_0_(cbx_4__7__1_top_grid_bottom_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_13__pin_f2a_i_0_(cbx_4__7__1_top_grid_bottom_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_14__pin_f2a_i_0_(cbx_4__7__1_top_grid_bottom_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_15__pin_f2a_i_0_(cbx_4__7__1_top_grid_bottom_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_16__pin_f2a_i_0_(cbx_4__7__1_top_grid_bottom_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_17__pin_f2a_i_0_(cbx_4__7__1_top_grid_bottom_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_18__pin_f2a_i_0_(cbx_4__7__1_top_grid_bottom_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_19__pin_f2a_i_0_(cbx_4__7__1_top_grid_bottom_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.ccff_tail(cbx_4__7__1_ccff_tail));

	cbx_7__1_ cbx_7__1_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chanx_left_in(sb_2__1__2_chanx_right_out[0:95]),
		.chanx_right_in(sb_7__1__0_chanx_left_out[0:95]),
		.ccff_head(sb_7__1__0_ccff_tail),
		.chanx_left_out(cbx_7__1__0_chanx_left_out[0:95]),
		.chanx_right_out(cbx_7__1__0_chanx_right_out[0:95]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_WDATA_A1_i_0_(cbx_7__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_WDATA_A1_i_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_WDATA_A1_i_1_(cbx_7__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_WDATA_A1_i_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_WDATA_A1_i_2_(cbx_7__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_WDATA_A1_i_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_WDATA_A1_i_3_(cbx_7__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_WDATA_A1_i_3_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_WDATA_A1_i_4_(cbx_7__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_WDATA_A1_i_4_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_WDATA_A1_i_5_(cbx_7__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_WDATA_A1_i_5_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_WDATA_A1_i_6_(cbx_7__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_WDATA_A1_i_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_6_(cbx_7__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_7_(cbx_7__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_7_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_8_(cbx_7__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_8_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_9_(cbx_7__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_9_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_10_(cbx_7__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_11_(cbx_7__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_11_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_12_(cbx_7__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_12_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_13_(cbx_7__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_13_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_14_(cbx_7__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_WDATA_B1_i_17_(cbx_7__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_WDATA_B1_i_17_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ADDR_B1_i_1_(cbx_7__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ADDR_B1_i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_f2a_i_0_(cbx_7__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_f2a_i_0_(cbx_7__1__0_bottom_grid_top_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_f2a_i_0_(cbx_7__1__0_bottom_grid_top_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_f2a_i_0_(cbx_7__1__0_bottom_grid_top_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_f2a_i_0_(cbx_7__1__0_bottom_grid_top_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_f2a_i_0_(cbx_7__1__0_bottom_grid_top_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_f2a_i_0_(cbx_7__1__0_bottom_grid_top_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_f2a_i_0_(cbx_7__1__0_bottom_grid_top_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_8__pin_f2a_i_0_(cbx_7__1__0_bottom_grid_top_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_9__pin_f2a_i_0_(cbx_7__1__0_bottom_grid_top_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_10__pin_f2a_i_0_(cbx_7__1__0_bottom_grid_top_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_11__pin_f2a_i_0_(cbx_7__1__0_bottom_grid_top_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_12__pin_f2a_i_0_(cbx_7__1__0_bottom_grid_top_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_13__pin_f2a_i_0_(cbx_7__1__0_bottom_grid_top_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_14__pin_f2a_i_0_(cbx_7__1__0_bottom_grid_top_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_15__pin_f2a_i_0_(cbx_7__1__0_bottom_grid_top_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_16__pin_f2a_i_0_(cbx_7__1__0_bottom_grid_top_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_17__pin_f2a_i_0_(cbx_7__1__0_bottom_grid_top_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_18__pin_f2a_i_0_(cbx_7__1__0_bottom_grid_top_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.bottom_grid_top_width_0_height_0_subtile_19__pin_f2a_i_0_(cbx_7__1__0_bottom_grid_top_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.ccff_tail(cbx_7__1__0_ccff_tail));

	cby_0__1_ cby_0__1_ (
		.chany_bottom_in(sb_0__0__0_chany_top_out[0:95]),
		.chany_top_in(sb_0__1__0_chany_bottom_out[0:95]),
		.chany_bottom_out(cby_0__1__0_chany_bottom_out[0:95]),
		.chany_top_out(cby_0__1__0_chany_top_out[0:95]));

	cby_0__1_ cby_0__2_ (
		.chany_bottom_in(sb_0__1__0_chany_top_out[0:95]),
		.chany_top_in(sb_0__1__1_chany_bottom_out[0:95]),
		.chany_bottom_out(cby_0__1__1_chany_bottom_out[0:95]),
		.chany_top_out(cby_0__1__1_chany_top_out[0:95]));

	cby_0__1_ cby_0__3_ (
		.chany_bottom_in(sb_0__1__1_chany_top_out[0:95]),
		.chany_top_in(sb_0__1__2_chany_bottom_out[0:95]),
		.chany_bottom_out(cby_0__1__2_chany_bottom_out[0:95]),
		.chany_top_out(cby_0__1__2_chany_top_out[0:95]));

	cby_0__1_ cby_0__4_ (
		.chany_bottom_in(sb_0__1__2_chany_top_out[0:95]),
		.chany_top_in(sb_0__1__3_chany_bottom_out[0:95]),
		.chany_bottom_out(cby_0__1__3_chany_bottom_out[0:95]),
		.chany_top_out(cby_0__1__3_chany_top_out[0:95]));

	cby_0__1_ cby_0__5_ (
		.chany_bottom_in(sb_0__1__3_chany_top_out[0:95]),
		.chany_top_in(sb_0__1__4_chany_bottom_out[0:95]),
		.chany_bottom_out(cby_0__1__4_chany_bottom_out[0:95]),
		.chany_top_out(cby_0__1__4_chany_top_out[0:95]));

	cby_0__1_ cby_0__6_ (
		.chany_bottom_in(sb_0__1__4_chany_top_out[0:95]),
		.chany_top_in(sb_0__1__5_chany_bottom_out[0:95]),
		.chany_bottom_out(cby_0__1__5_chany_bottom_out[0:95]),
		.chany_top_out(cby_0__1__5_chany_top_out[0:95]));

	cby_0__1_ cby_0__7_ (
		.chany_bottom_in(sb_0__1__5_chany_top_out[0:95]),
		.chany_top_in(sb_0__1__6_chany_bottom_out[0:95]),
		.chany_bottom_out(cby_0__1__6_chany_bottom_out[0:95]),
		.chany_top_out(cby_0__1__6_chany_top_out[0:95]));

	cby_0__1_ cby_0__8_ (
		.chany_bottom_in(sb_0__1__6_chany_top_out[0:95]),
		.chany_top_in(sb_0__8__0_chany_bottom_out[0:95]),
		.chany_bottom_out(cby_0__1__7_chany_bottom_out[0:95]),
		.chany_top_out(cby_0__1__7_chany_top_out[0:95]));

	cby_0__1_ cby_2__1_ (
		.chany_bottom_in(sb_2__0__0_chany_top_out[0:95]),
		.chany_top_in(sb_2__1__0_chany_bottom_out[0:95]),
		.chany_bottom_out(cby_0__1__8_chany_bottom_out[0:95]),
		.chany_top_out(cby_0__1__8_chany_top_out[0:95]));

	cby_0__1_ cby_2__8_ (
		.chany_bottom_in(sb_2__7__0_chany_top_out[0:95]),
		.chany_top_in(sb_2__8__0_chany_bottom_out[0:95]),
		.chany_bottom_out(cby_0__1__9_chany_bottom_out[0:95]),
		.chany_top_out(cby_0__1__9_chany_top_out[0:95]));

	cby_0__1_ cby_3__1_ (
		.chany_bottom_in(sb_2__0__1_chany_top_out[0:95]),
		.chany_top_in(sb_3__1__0_chany_bottom_out[0:95]),
		.chany_bottom_out(cby_0__1__10_chany_bottom_out[0:95]),
		.chany_top_out(cby_0__1__10_chany_top_out[0:95]));

	cby_0__1_ cby_3__8_ (
		.chany_bottom_in(sb_3__7__0_chany_top_out[0:95]),
		.chany_top_in(sb_2__8__1_chany_bottom_out[0:95]),
		.chany_bottom_out(cby_0__1__11_chany_bottom_out[0:95]),
		.chany_top_out(cby_0__1__11_chany_top_out[0:95]));

	cby_0__1_ cby_4__1_ (
		.chany_bottom_in(sb_2__0__2_chany_top_out[0:95]),
		.chany_top_in(sb_4__1__0_chany_bottom_out[0:95]),
		.chany_bottom_out(cby_0__1__12_chany_bottom_out[0:95]),
		.chany_top_out(cby_0__1__12_chany_top_out[0:95]));

	cby_0__1_ cby_4__8_ (
		.chany_bottom_in(sb_4__7__0_chany_top_out[0:95]),
		.chany_top_in(sb_2__8__2_chany_bottom_out[0:95]),
		.chany_bottom_out(cby_0__1__13_chany_bottom_out[0:95]),
		.chany_top_out(cby_0__1__13_chany_top_out[0:95]));

	cby_0__1_ cby_5__1_ (
		.chany_bottom_in(sb_2__0__3_chany_top_out[0:95]),
		.chany_top_in(sb_2__1__1_chany_bottom_out[0:95]),
		.chany_bottom_out(cby_0__1__14_chany_bottom_out[0:95]),
		.chany_top_out(cby_0__1__14_chany_top_out[0:95]));

	cby_0__1_ cby_5__8_ (
		.chany_bottom_in(sb_2__7__1_chany_top_out[0:95]),
		.chany_top_in(sb_2__8__3_chany_bottom_out[0:95]),
		.chany_bottom_out(cby_0__1__15_chany_bottom_out[0:95]),
		.chany_top_out(cby_0__1__15_chany_top_out[0:95]));

	cby_0__1_ cby_6__1_ (
		.chany_bottom_in(sb_2__0__4_chany_top_out[0:95]),
		.chany_top_in(sb_2__1__2_chany_bottom_out[0:95]),
		.chany_bottom_out(cby_0__1__16_chany_bottom_out[0:95]),
		.chany_top_out(cby_0__1__16_chany_top_out[0:95]));

	cby_0__1_ cby_6__8_ (
		.chany_bottom_in(sb_3__7__1_chany_top_out[0:95]),
		.chany_top_in(sb_2__8__4_chany_bottom_out[0:95]),
		.chany_bottom_out(cby_0__1__17_chany_bottom_out[0:95]),
		.chany_top_out(cby_0__1__17_chany_top_out[0:95]));

	cby_0__1_ cby_7__1_ (
		.chany_bottom_in(sb_2__0__5_chany_top_out[0:95]),
		.chany_top_in(sb_7__1__0_chany_bottom_out[0:95]),
		.chany_bottom_out(cby_0__1__18_chany_bottom_out[0:95]),
		.chany_top_out(cby_0__1__18_chany_top_out[0:95]));

	cby_0__1_ cby_7__8_ (
		.chany_bottom_in(sb_7__7__0_chany_top_out[0:95]),
		.chany_top_in(sb_2__8__5_chany_bottom_out[0:95]),
		.chany_bottom_out(cby_0__1__19_chany_bottom_out[0:95]),
		.chany_top_out(cby_0__1__19_chany_top_out[0:95]));

	cby_0__1_ cby_8__1_ (
		.chany_bottom_in(sb_2__0__6_chany_top_out[0:95]),
		.chany_top_in(sb_2__1__3_chany_bottom_out[0:95]),
		.chany_bottom_out(cby_0__1__20_chany_bottom_out[0:95]),
		.chany_top_out(cby_0__1__20_chany_top_out[0:95]));

	cby_0__1_ cby_8__8_ (
		.chany_bottom_in(sb_2__7__2_chany_top_out[0:95]),
		.chany_top_in(sb_2__8__6_chany_bottom_out[0:95]),
		.chany_bottom_out(cby_0__1__21_chany_bottom_out[0:95]),
		.chany_top_out(cby_0__1__21_chany_top_out[0:95]));

	cby_0__1_ cby_10__1_ (
		.chany_bottom_in(sb_10__0__0_chany_top_out[0:95]),
		.chany_top_in(sb_10__1__0_chany_bottom_out[0:95]),
		.chany_bottom_out(cby_0__1__22_chany_bottom_out[0:95]),
		.chany_top_out(cby_0__1__22_chany_top_out[0:95]));

	cby_0__1_ cby_10__2_ (
		.chany_bottom_in(sb_10__1__0_chany_top_out[0:95]),
		.chany_top_in(sb_10__1__1_chany_bottom_out[0:95]),
		.chany_bottom_out(cby_0__1__23_chany_bottom_out[0:95]),
		.chany_top_out(cby_0__1__23_chany_top_out[0:95]));

	cby_0__1_ cby_10__3_ (
		.chany_bottom_in(sb_10__1__1_chany_top_out[0:95]),
		.chany_top_in(sb_10__1__2_chany_bottom_out[0:95]),
		.chany_bottom_out(cby_0__1__24_chany_bottom_out[0:95]),
		.chany_top_out(cby_0__1__24_chany_top_out[0:95]));

	cby_0__1_ cby_10__4_ (
		.chany_bottom_in(sb_10__1__2_chany_top_out[0:95]),
		.chany_top_in(sb_10__1__3_chany_bottom_out[0:95]),
		.chany_bottom_out(cby_0__1__25_chany_bottom_out[0:95]),
		.chany_top_out(cby_0__1__25_chany_top_out[0:95]));

	cby_0__1_ cby_10__5_ (
		.chany_bottom_in(sb_10__1__3_chany_top_out[0:95]),
		.chany_top_in(sb_10__1__4_chany_bottom_out[0:95]),
		.chany_bottom_out(cby_0__1__26_chany_bottom_out[0:95]),
		.chany_top_out(cby_0__1__26_chany_top_out[0:95]));

	cby_0__1_ cby_10__6_ (
		.chany_bottom_in(sb_10__1__4_chany_top_out[0:95]),
		.chany_top_in(sb_10__1__5_chany_bottom_out[0:95]),
		.chany_bottom_out(cby_0__1__27_chany_bottom_out[0:95]),
		.chany_top_out(cby_0__1__27_chany_top_out[0:95]));

	cby_0__1_ cby_10__7_ (
		.chany_bottom_in(sb_10__1__5_chany_top_out[0:95]),
		.chany_top_in(sb_10__1__6_chany_bottom_out[0:95]),
		.chany_bottom_out(cby_0__1__28_chany_bottom_out[0:95]),
		.chany_top_out(cby_0__1__28_chany_top_out[0:95]));

	cby_0__1_ cby_10__8_ (
		.chany_bottom_in(sb_10__1__6_chany_top_out[0:95]),
		.chany_top_in(sb_10__8__0_chany_bottom_out[0:95]),
		.chany_bottom_out(cby_0__1__29_chany_bottom_out[0:95]),
		.chany_top_out(cby_0__1__29_chany_top_out[0:95]));

	cby_1__1_ cby_1__1_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_bottom_in(sb_1__0__0_chany_top_out[0:95]),
		.chany_top_in(sb_1__1__0_chany_bottom_out[0:95]),
		.ccff_head(sb_1__0__0_ccff_tail),
		.chany_bottom_out(cby_1__1__0_chany_bottom_out[0:95]),
		.chany_top_out(cby_1__1__0_chany_top_out[0:95]),
		.left_grid_right_width_0_height_0_subtile_0__pin_f2a_i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_f2a_i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_f2a_i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_f2a_i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_f2a_i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_f2a_i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_f2a_i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_f2a_i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_8__pin_f2a_i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_9__pin_f2a_i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_10__pin_f2a_i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_11__pin_f2a_i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_12__pin_f2a_i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_13__pin_f2a_i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_14__pin_f2a_i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_15__pin_f2a_i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_16__pin_f2a_i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_17__pin_f2a_i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_18__pin_f2a_i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_19__pin_f2a_i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.ccff_tail(cby_1__1__0_ccff_tail));

	cby_1__1_ cby_1__2_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_bottom_in(sb_1__1__0_chany_top_out[0:95]),
		.chany_top_in(sb_1__2__0_chany_bottom_out[0:95]),
		.ccff_head(sb_1__1__0_ccff_tail),
		.chany_bottom_out(cby_1__1__1_chany_bottom_out[0:95]),
		.chany_top_out(cby_1__1__1_chany_top_out[0:95]),
		.left_grid_right_width_0_height_0_subtile_0__pin_f2a_i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_f2a_i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_f2a_i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_f2a_i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_f2a_i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_f2a_i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_f2a_i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_f2a_i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_8__pin_f2a_i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_9__pin_f2a_i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_10__pin_f2a_i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_11__pin_f2a_i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_12__pin_f2a_i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_13__pin_f2a_i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_14__pin_f2a_i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_15__pin_f2a_i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_16__pin_f2a_i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_17__pin_f2a_i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_18__pin_f2a_i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_19__pin_f2a_i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.ccff_tail(cby_1__1__1_ccff_tail));

	cby_1__1_ cby_1__3_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_bottom_in(sb_1__2__0_chany_top_out[0:95]),
		.chany_top_in(sb_1__2__1_chany_bottom_out[0:95]),
		.ccff_head(sb_1__2__0_ccff_tail),
		.chany_bottom_out(cby_1__1__2_chany_bottom_out[0:95]),
		.chany_top_out(cby_1__1__2_chany_top_out[0:95]),
		.left_grid_right_width_0_height_0_subtile_0__pin_f2a_i_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_f2a_i_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_f2a_i_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_f2a_i_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_f2a_i_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_f2a_i_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_f2a_i_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_f2a_i_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_8__pin_f2a_i_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_9__pin_f2a_i_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_10__pin_f2a_i_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_11__pin_f2a_i_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_12__pin_f2a_i_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_13__pin_f2a_i_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_14__pin_f2a_i_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_15__pin_f2a_i_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_16__pin_f2a_i_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_17__pin_f2a_i_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_18__pin_f2a_i_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_19__pin_f2a_i_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.ccff_tail(cby_1__1__2_ccff_tail));

	cby_1__1_ cby_1__4_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_bottom_in(sb_1__2__1_chany_top_out[0:95]),
		.chany_top_in(sb_1__2__2_chany_bottom_out[0:95]),
		.ccff_head(sb_1__2__1_ccff_tail),
		.chany_bottom_out(cby_1__1__3_chany_bottom_out[0:95]),
		.chany_top_out(cby_1__1__3_chany_top_out[0:95]),
		.left_grid_right_width_0_height_0_subtile_0__pin_f2a_i_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_f2a_i_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_f2a_i_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_f2a_i_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_f2a_i_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_f2a_i_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_f2a_i_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_f2a_i_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_8__pin_f2a_i_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_9__pin_f2a_i_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_10__pin_f2a_i_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_11__pin_f2a_i_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_12__pin_f2a_i_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_13__pin_f2a_i_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_14__pin_f2a_i_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_15__pin_f2a_i_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_16__pin_f2a_i_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_17__pin_f2a_i_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_18__pin_f2a_i_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_19__pin_f2a_i_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.ccff_tail(cby_1__1__3_ccff_tail));

	cby_1__1_ cby_1__5_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_bottom_in(sb_1__2__2_chany_top_out[0:95]),
		.chany_top_in(sb_1__2__3_chany_bottom_out[0:95]),
		.ccff_head(sb_1__2__2_ccff_tail),
		.chany_bottom_out(cby_1__1__4_chany_bottom_out[0:95]),
		.chany_top_out(cby_1__1__4_chany_top_out[0:95]),
		.left_grid_right_width_0_height_0_subtile_0__pin_f2a_i_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_f2a_i_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_f2a_i_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_f2a_i_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_f2a_i_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_f2a_i_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_f2a_i_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_f2a_i_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_8__pin_f2a_i_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_9__pin_f2a_i_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_10__pin_f2a_i_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_11__pin_f2a_i_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_12__pin_f2a_i_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_13__pin_f2a_i_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_14__pin_f2a_i_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_15__pin_f2a_i_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_16__pin_f2a_i_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_17__pin_f2a_i_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_18__pin_f2a_i_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_19__pin_f2a_i_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.ccff_tail(cby_1__1__4_ccff_tail));

	cby_1__1_ cby_1__6_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_bottom_in(sb_1__2__3_chany_top_out[0:95]),
		.chany_top_in(sb_1__2__4_chany_bottom_out[0:95]),
		.ccff_head(sb_1__2__3_ccff_tail),
		.chany_bottom_out(cby_1__1__5_chany_bottom_out[0:95]),
		.chany_top_out(cby_1__1__5_chany_top_out[0:95]),
		.left_grid_right_width_0_height_0_subtile_0__pin_f2a_i_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_f2a_i_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_f2a_i_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_f2a_i_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_f2a_i_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_f2a_i_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_f2a_i_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_f2a_i_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_8__pin_f2a_i_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_9__pin_f2a_i_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_10__pin_f2a_i_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_11__pin_f2a_i_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_12__pin_f2a_i_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_13__pin_f2a_i_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_14__pin_f2a_i_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_15__pin_f2a_i_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_16__pin_f2a_i_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_17__pin_f2a_i_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_18__pin_f2a_i_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_19__pin_f2a_i_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.ccff_tail(cby_1__1__5_ccff_tail));

	cby_1__1_ cby_1__7_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_bottom_in(sb_1__2__4_chany_top_out[0:95]),
		.chany_top_in(sb_1__7__0_chany_bottom_out[0:95]),
		.ccff_head(sb_1__2__4_ccff_tail),
		.chany_bottom_out(cby_1__1__6_chany_bottom_out[0:95]),
		.chany_top_out(cby_1__1__6_chany_top_out[0:95]),
		.left_grid_right_width_0_height_0_subtile_0__pin_f2a_i_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_f2a_i_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_f2a_i_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_f2a_i_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_f2a_i_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_f2a_i_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_f2a_i_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_f2a_i_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_8__pin_f2a_i_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_9__pin_f2a_i_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_10__pin_f2a_i_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_11__pin_f2a_i_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_12__pin_f2a_i_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_13__pin_f2a_i_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_14__pin_f2a_i_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_15__pin_f2a_i_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_16__pin_f2a_i_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_17__pin_f2a_i_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_18__pin_f2a_i_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_19__pin_f2a_i_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.ccff_tail(cby_1__1__6_ccff_tail));

	cby_1__1_ cby_1__8_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_bottom_in(sb_1__7__0_chany_top_out[0:95]),
		.chany_top_in(sb_1__8__0_chany_bottom_out[0:95]),
		.ccff_head(sb_1__7__0_ccff_tail),
		.chany_bottom_out(cby_1__1__7_chany_bottom_out[0:95]),
		.chany_top_out(cby_1__1__7_chany_top_out[0:95]),
		.left_grid_right_width_0_height_0_subtile_0__pin_f2a_i_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_f2a_i_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_f2a_i_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_f2a_i_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_f2a_i_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_f2a_i_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_f2a_i_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_f2a_i_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_8__pin_f2a_i_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_9__pin_f2a_i_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_10__pin_f2a_i_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_11__pin_f2a_i_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_12__pin_f2a_i_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_13__pin_f2a_i_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_14__pin_f2a_i_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_15__pin_f2a_i_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_16__pin_f2a_i_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_17__pin_f2a_i_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_18__pin_f2a_i_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_19__pin_f2a_i_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.ccff_tail(cby_1__1__7_ccff_tail));

	cby_2__2_ cby_2__2_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_bottom_in(sb_2__1__0_chany_top_out[0:95]),
		.chany_top_in(sb_2__2__0_chany_bottom_out[0:95]),
		.ccff_head(cbx_2__1__0_ccff_tail),
		.chany_bottom_out(cby_2__2__0_chany_bottom_out[0:95]),
		.chany_top_out(cby_2__2__0_chany_top_out[0:95]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__0_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__0_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__0_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__0_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__0_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__0_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.ccff_tail(cby_2__2__0_ccff_tail));

	cby_2__2_ cby_2__3_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_bottom_in(sb_2__2__0_chany_top_out[0:95]),
		.chany_top_in(sb_2__2__1_chany_bottom_out[0:95]),
		.ccff_head(cbx_2__2__0_ccff_tail),
		.chany_bottom_out(cby_2__2__1_chany_bottom_out[0:95]),
		.chany_top_out(cby_2__2__1_chany_top_out[0:95]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__1_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__1_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__1_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__1_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__1_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__1_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.ccff_tail(cby_2__2__1_ccff_tail));

	cby_2__2_ cby_2__4_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_bottom_in(sb_2__2__1_chany_top_out[0:95]),
		.chany_top_in(sb_2__2__2_chany_bottom_out[0:95]),
		.ccff_head(ccff_head[5]),
		.chany_bottom_out(cby_2__2__2_chany_bottom_out[0:95]),
		.chany_top_out(cby_2__2__2_chany_top_out[0:95]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__2_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__2_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__2_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__2_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__2_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__2_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.ccff_tail(cby_2__2__2_ccff_tail));

	cby_2__2_ cby_2__5_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_bottom_in(sb_2__2__2_chany_top_out[0:95]),
		.chany_top_in(sb_2__2__3_chany_bottom_out[0:95]),
		.ccff_head(cbx_2__2__2_ccff_tail),
		.chany_bottom_out(cby_2__2__3_chany_bottom_out[0:95]),
		.chany_top_out(cby_2__2__3_chany_top_out[0:95]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__3_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__3_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__3_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__3_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__3_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__3_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.ccff_tail(cby_2__2__3_ccff_tail));

	cby_2__2_ cby_2__6_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_bottom_in(sb_2__2__3_chany_top_out[0:95]),
		.chany_top_in(sb_2__2__4_chany_bottom_out[0:95]),
		.ccff_head(cbx_2__2__3_ccff_tail),
		.chany_bottom_out(cby_2__2__4_chany_bottom_out[0:95]),
		.chany_top_out(cby_2__2__4_chany_top_out[0:95]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__4_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__4_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__4_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__4_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__4_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__4_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.ccff_tail(cby_2__2__4_ccff_tail));

	cby_2__2_ cby_2__7_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_bottom_in(sb_2__2__4_chany_top_out[0:95]),
		.chany_top_in(sb_2__7__0_chany_bottom_out[0:95]),
		.ccff_head(cbx_2__2__4_ccff_tail),
		.chany_bottom_out(cby_2__2__5_chany_bottom_out[0:95]),
		.chany_top_out(cby_2__2__5_chany_top_out[0:95]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__5_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__5_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__5_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__5_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__5_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__5_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.ccff_tail(cby_2__2__5_ccff_tail));

	cby_2__2_ cby_3__2_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_bottom_in(sb_3__1__0_chany_top_out[0:95]),
		.chany_top_in(sb_3__2__0_chany_bottom_out[0:95]),
		.ccff_head(cbx_2__1__1_ccff_tail),
		.chany_bottom_out(cby_2__2__6_chany_bottom_out[0:95]),
		.chany_top_out(cby_2__2__6_chany_top_out[0:95]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__6_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__6_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__6_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__6_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__6_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__6_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__6_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.ccff_tail(cby_2__2__6_ccff_tail));

	cby_2__2_ cby_3__3_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_bottom_in(sb_3__2__0_chany_top_out[0:95]),
		.chany_top_in(sb_3__2__1_chany_bottom_out[0:95]),
		.ccff_head(cbx_2__2__5_ccff_tail),
		.chany_bottom_out(cby_2__2__7_chany_bottom_out[0:95]),
		.chany_top_out(cby_2__2__7_chany_top_out[0:95]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__7_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__7_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__7_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__7_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__7_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__7_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__7_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.ccff_tail(cby_2__2__7_ccff_tail));

	cby_2__2_ cby_3__4_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_bottom_in(sb_3__2__1_chany_top_out[0:95]),
		.chany_top_in(sb_3__4__0_chany_bottom_out[0:95]),
		.ccff_head(cbx_2__2__6_ccff_tail),
		.chany_bottom_out(cby_2__2__8_chany_bottom_out[0:95]),
		.chany_top_out(cby_2__2__8_chany_top_out[0:95]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__8_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__8_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__8_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__8_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__8_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__8_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__8_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.ccff_tail(cby_2__2__8_ccff_tail));

	cby_2__2_ cby_3__5_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_bottom_in(sb_3__4__0_chany_top_out[0:95]),
		.chany_top_in(sb_3__2__2_chany_bottom_out[0:95]),
		.ccff_head(cbx_2__2__7_ccff_tail),
		.chany_bottom_out(cby_2__2__9_chany_bottom_out[0:95]),
		.chany_top_out(cby_2__2__9_chany_top_out[0:95]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__9_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__9_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__9_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__9_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__9_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__9_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__9_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.ccff_tail(cby_2__2__9_ccff_tail));

	cby_2__2_ cby_3__6_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_bottom_in(sb_3__2__2_chany_top_out[0:95]),
		.chany_top_in(sb_3__2__3_chany_bottom_out[0:95]),
		.ccff_head(cbx_2__2__8_ccff_tail),
		.chany_bottom_out(cby_2__2__10_chany_bottom_out[0:95]),
		.chany_top_out(cby_2__2__10_chany_top_out[0:95]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__10_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__10_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__10_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__10_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__10_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__10_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__10_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.ccff_tail(cby_2__2__10_ccff_tail));

	cby_2__2_ cby_3__7_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_bottom_in(sb_3__2__3_chany_top_out[0:95]),
		.chany_top_in(sb_3__7__0_chany_bottom_out[0:95]),
		.ccff_head(cbx_2__2__9_ccff_tail),
		.chany_bottom_out(cby_2__2__11_chany_bottom_out[0:95]),
		.chany_top_out(cby_2__2__11_chany_top_out[0:95]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__11_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__11_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__11_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__11_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__11_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__11_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__11_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.ccff_tail(cby_2__2__11_ccff_tail));

	cby_2__2_ cby_5__2_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_bottom_in(sb_2__1__1_chany_top_out[0:95]),
		.chany_top_in(sb_2__2__5_chany_bottom_out[0:95]),
		.ccff_head(cbx_2__1__2_ccff_tail),
		.chany_bottom_out(cby_2__2__12_chany_bottom_out[0:95]),
		.chany_top_out(cby_2__2__12_chany_top_out[0:95]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__12_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__12_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__12_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__12_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__12_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__12_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__12_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.ccff_tail(cby_2__2__12_ccff_tail));

	cby_2__2_ cby_5__3_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_bottom_in(sb_2__2__5_chany_top_out[0:95]),
		.chany_top_in(sb_2__2__6_chany_bottom_out[0:95]),
		.ccff_head(cbx_2__2__10_ccff_tail),
		.chany_bottom_out(cby_2__2__13_chany_bottom_out[0:95]),
		.chany_top_out(cby_2__2__13_chany_top_out[0:95]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__13_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__13_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__13_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__13_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__13_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__13_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__13_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.ccff_tail(cby_2__2__13_ccff_tail));

	cby_2__2_ cby_5__4_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_bottom_in(sb_2__2__6_chany_top_out[0:95]),
		.chany_top_in(sb_2__2__7_chany_bottom_out[0:95]),
		.ccff_head(cbx_2__2__11_ccff_tail),
		.chany_bottom_out(cby_2__2__14_chany_bottom_out[0:95]),
		.chany_top_out(cby_2__2__14_chany_top_out[0:95]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__14_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__14_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__14_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__14_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__14_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__14_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__14_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.ccff_tail(cby_2__2__14_ccff_tail));

	cby_2__2_ cby_5__5_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_bottom_in(sb_2__2__7_chany_top_out[0:95]),
		.chany_top_in(sb_2__2__8_chany_bottom_out[0:95]),
		.ccff_head(cbx_2__2__12_ccff_tail),
		.chany_bottom_out(cby_2__2__15_chany_bottom_out[0:95]),
		.chany_top_out(cby_2__2__15_chany_top_out[0:95]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__15_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__15_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__15_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__15_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__15_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__15_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__15_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.ccff_tail(cby_2__2__15_ccff_tail));

	cby_2__2_ cby_5__6_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_bottom_in(sb_2__2__8_chany_top_out[0:95]),
		.chany_top_in(sb_2__2__9_chany_bottom_out[0:95]),
		.ccff_head(cbx_2__2__13_ccff_tail),
		.chany_bottom_out(cby_2__2__16_chany_bottom_out[0:95]),
		.chany_top_out(cby_2__2__16_chany_top_out[0:95]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__16_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__16_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__16_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__16_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__16_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__16_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__16_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.ccff_tail(cby_2__2__16_ccff_tail));

	cby_2__2_ cby_5__7_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_bottom_in(sb_2__2__9_chany_top_out[0:95]),
		.chany_top_in(sb_2__7__1_chany_bottom_out[0:95]),
		.ccff_head(cbx_2__2__14_ccff_tail),
		.chany_bottom_out(cby_2__2__17_chany_bottom_out[0:95]),
		.chany_top_out(cby_2__2__17_chany_top_out[0:95]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__17_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__17_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__17_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__17_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__17_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__17_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__17_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.ccff_tail(cby_2__2__17_ccff_tail));

	cby_2__2_ cby_6__2_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_bottom_in(sb_2__1__2_chany_top_out[0:95]),
		.chany_top_in(sb_3__2__4_chany_bottom_out[0:95]),
		.ccff_head(cbx_2__1__3_ccff_tail),
		.chany_bottom_out(cby_2__2__18_chany_bottom_out[0:95]),
		.chany_top_out(cby_2__2__18_chany_top_out[0:95]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__18_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__18_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__18_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__18_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__18_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__18_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__18_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__18_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__18_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__18_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__18_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__18_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__18_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__18_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__18_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__18_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__18_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__18_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__18_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__18_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__18_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__18_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__18_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__18_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__18_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__18_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.ccff_tail(ccff_tail[1]));

	cby_2__2_ cby_6__3_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_bottom_in(sb_3__2__4_chany_top_out[0:95]),
		.chany_top_in(sb_3__2__5_chany_bottom_out[0:95]),
		.ccff_head(cbx_2__2__15_ccff_tail),
		.chany_bottom_out(cby_2__2__19_chany_bottom_out[0:95]),
		.chany_top_out(cby_2__2__19_chany_top_out[0:95]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__19_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__19_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__19_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__19_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__19_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__19_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__19_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__19_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__19_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__19_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__19_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__19_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__19_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__19_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__19_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__19_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__19_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__19_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__19_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__19_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__19_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__19_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__19_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__19_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__19_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__19_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.ccff_tail(cby_2__2__19_ccff_tail));

	cby_2__2_ cby_6__4_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_bottom_in(sb_3__2__5_chany_top_out[0:95]),
		.chany_top_in(sb_3__2__6_chany_bottom_out[0:95]),
		.ccff_head(cbx_2__2__16_ccff_tail),
		.chany_bottom_out(cby_2__2__20_chany_bottom_out[0:95]),
		.chany_top_out(cby_2__2__20_chany_top_out[0:95]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__20_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__20_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__20_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__20_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__20_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__20_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__20_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__20_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__20_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__20_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__20_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__20_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__20_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__20_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__20_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__20_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__20_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__20_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__20_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__20_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__20_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__20_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__20_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__20_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__20_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__20_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.ccff_tail(cby_2__2__20_ccff_tail));

	cby_2__2_ cby_6__5_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_bottom_in(sb_3__2__6_chany_top_out[0:95]),
		.chany_top_in(sb_3__2__7_chany_bottom_out[0:95]),
		.ccff_head(cbx_2__2__17_ccff_tail),
		.chany_bottom_out(cby_2__2__21_chany_bottom_out[0:95]),
		.chany_top_out(cby_2__2__21_chany_top_out[0:95]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__21_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__21_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__21_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__21_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__21_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__21_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__21_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__21_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__21_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__21_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__21_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__21_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__21_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__21_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__21_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__21_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__21_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__21_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__21_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__21_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__21_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__21_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__21_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__21_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__21_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__21_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.ccff_tail(ccff_tail[5]));

	cby_2__2_ cby_6__6_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_bottom_in(sb_3__2__7_chany_top_out[0:95]),
		.chany_top_in(sb_3__2__8_chany_bottom_out[0:95]),
		.ccff_head(ccff_head[7]),
		.chany_bottom_out(cby_2__2__22_chany_bottom_out[0:95]),
		.chany_top_out(cby_2__2__22_chany_top_out[0:95]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__22_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__22_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__22_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__22_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__22_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__22_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__22_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__22_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__22_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__22_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__22_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__22_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__22_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__22_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__22_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__22_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__22_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__22_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__22_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__22_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__22_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__22_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__22_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__22_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__22_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__22_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.ccff_tail(cby_2__2__22_ccff_tail));

	cby_2__2_ cby_6__7_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_bottom_in(sb_3__2__8_chany_top_out[0:95]),
		.chany_top_in(sb_3__7__1_chany_bottom_out[0:95]),
		.ccff_head(cbx_2__2__19_ccff_tail),
		.chany_bottom_out(cby_2__2__23_chany_bottom_out[0:95]),
		.chany_top_out(cby_2__2__23_chany_top_out[0:95]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__23_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__23_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__23_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__23_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__23_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__23_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__23_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__23_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__23_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__23_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__23_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__23_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__23_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__23_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__23_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__23_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__23_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__23_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__23_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__23_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__23_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__23_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__23_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__23_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__23_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__23_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.ccff_tail(cby_2__2__23_ccff_tail));

	cby_2__2_ cby_8__2_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_bottom_in(sb_2__1__3_chany_top_out[0:95]),
		.chany_top_in(sb_2__2__10_chany_bottom_out[0:95]),
		.ccff_head(cbx_2__1__4_ccff_tail),
		.chany_bottom_out(cby_2__2__24_chany_bottom_out[0:95]),
		.chany_top_out(cby_2__2__24_chany_top_out[0:95]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__24_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__24_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__24_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__24_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__24_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__24_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__24_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__24_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__24_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__24_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__24_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__24_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__24_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__24_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__24_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__24_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__24_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__24_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__24_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__24_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__24_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__24_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__24_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__24_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__24_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__24_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.ccff_tail(cby_2__2__24_ccff_tail));

	cby_2__2_ cby_8__3_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_bottom_in(sb_2__2__10_chany_top_out[0:95]),
		.chany_top_in(sb_2__2__11_chany_bottom_out[0:95]),
		.ccff_head(cbx_2__2__20_ccff_tail),
		.chany_bottom_out(cby_2__2__25_chany_bottom_out[0:95]),
		.chany_top_out(cby_2__2__25_chany_top_out[0:95]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__25_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__25_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__25_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__25_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__25_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__25_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__25_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__25_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__25_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__25_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__25_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__25_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__25_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__25_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__25_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__25_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__25_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__25_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__25_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__25_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__25_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__25_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__25_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__25_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__25_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__25_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.ccff_tail(cby_2__2__25_ccff_tail));

	cby_2__2_ cby_8__4_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_bottom_in(sb_2__2__11_chany_top_out[0:95]),
		.chany_top_in(sb_2__2__12_chany_bottom_out[0:95]),
		.ccff_head(cbx_2__2__21_ccff_tail),
		.chany_bottom_out(cby_2__2__26_chany_bottom_out[0:95]),
		.chany_top_out(cby_2__2__26_chany_top_out[0:95]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__26_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__26_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__26_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__26_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__26_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__26_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__26_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__26_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__26_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__26_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__26_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__26_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__26_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__26_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__26_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__26_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__26_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__26_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__26_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__26_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__26_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__26_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__26_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__26_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__26_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__26_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.ccff_tail(cby_2__2__26_ccff_tail));

	cby_2__2_ cby_8__5_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_bottom_in(sb_2__2__12_chany_top_out[0:95]),
		.chany_top_in(sb_2__2__13_chany_bottom_out[0:95]),
		.ccff_head(cbx_2__2__22_ccff_tail),
		.chany_bottom_out(cby_2__2__27_chany_bottom_out[0:95]),
		.chany_top_out(cby_2__2__27_chany_top_out[0:95]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__27_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__27_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__27_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__27_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__27_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__27_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__27_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__27_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__27_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__27_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__27_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__27_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__27_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__27_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__27_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__27_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__27_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__27_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__27_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__27_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__27_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__27_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__27_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__27_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__27_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__27_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.ccff_tail(cby_2__2__27_ccff_tail));

	cby_2__2_ cby_8__6_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_bottom_in(sb_2__2__13_chany_top_out[0:95]),
		.chany_top_in(sb_2__2__14_chany_bottom_out[0:95]),
		.ccff_head(cbx_2__2__23_ccff_tail),
		.chany_bottom_out(cby_2__2__28_chany_bottom_out[0:95]),
		.chany_top_out(cby_2__2__28_chany_top_out[0:95]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__28_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__28_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__28_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__28_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__28_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__28_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__28_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__28_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__28_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__28_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__28_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__28_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__28_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__28_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__28_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__28_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__28_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__28_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__28_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__28_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__28_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__28_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__28_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__28_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__28_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__28_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.ccff_tail(cby_2__2__28_ccff_tail));

	cby_2__2_ cby_8__7_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_bottom_in(sb_2__2__14_chany_top_out[0:95]),
		.chany_top_in(sb_2__7__2_chany_bottom_out[0:95]),
		.ccff_head(cbx_2__2__24_ccff_tail),
		.chany_bottom_out(cby_2__2__29_chany_bottom_out[0:95]),
		.chany_top_out(cby_2__2__29_chany_top_out[0:95]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_0_(cby_2__2__29_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_1_(cby_2__2__29_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_2_(cby_2__2__29_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_3_(cby_2__2__29_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_4_(cby_2__2__29_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_5_(cby_2__2__29_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_6_(cby_2__2__29_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_7_(cby_2__2__29_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_8_(cby_2__2__29_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_9_(cby_2__2__29_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_0_(cby_2__2__29_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_1_(cby_2__2__29_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_2_(cby_2__2__29_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_3_(cby_2__2__29_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_4_(cby_2__2__29_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_5_(cby_2__2__29_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_6_(cby_2__2__29_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_7_(cby_2__2__29_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_8_(cby_2__2__29_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_9_(cby_2__2__29_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_0_(cby_2__2__29_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_1_(cby_2__2__29_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_2_(cby_2__2__29_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_3_(cby_2__2__29_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_4_(cby_2__2__29_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_5_(cby_2__2__29_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.ccff_tail(cby_2__2__29_ccff_tail));

	cby_4__2_ cby_4__2_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_bottom_in(sb_4__1__0_chany_top_out[0:95]),
		.chany_top_in(sb_4__2__0_chany_bottom_out[0:95]),
		.ccff_head(cbx_4__1__0_ccff_tail),
		.chany_bottom_out(cby_4__2__0_chany_bottom_out[0:95]),
		.chany_top_out(cby_4__2__0_chany_top_out[0:95]),
		.left_grid_right_width_0_height_0_subtile_0__pin_a_i_2_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_a_i_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_a_i_3_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_a_i_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_a_i_4_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_a_i_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_a_i_5_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_a_i_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_a_i_6_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_a_i_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_a_i_7_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_a_i_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_acc_fir_i_1_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_acc_fir_i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_acc_fir_i_2_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_acc_fir_i_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_b_i_0_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_b_i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_b_i_1_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_b_i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_b_i_2_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_b_i_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_b_i_3_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_b_i_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_b_i_4_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_b_i_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_b_i_5_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_b_i_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_unsigned_a_0_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_unsigned_a_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_round_0_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_round_0_),
		.ccff_tail(cby_4__2__0_ccff_tail));

	cby_4__2_ cby_4__5_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_bottom_in(sb_4__4__0_chany_top_out[0:95]),
		.chany_top_in(sb_4__2__1_chany_bottom_out[0:95]),
		.ccff_head(cbx_4__4__0_ccff_tail),
		.chany_bottom_out(cby_4__2__1_chany_bottom_out[0:95]),
		.chany_top_out(cby_4__2__1_chany_top_out[0:95]),
		.left_grid_right_width_0_height_0_subtile_0__pin_a_i_2_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_a_i_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_a_i_3_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_a_i_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_a_i_4_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_a_i_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_a_i_5_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_a_i_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_a_i_6_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_a_i_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_a_i_7_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_a_i_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_acc_fir_i_1_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_acc_fir_i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_acc_fir_i_2_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_acc_fir_i_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_b_i_0_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_b_i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_b_i_1_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_b_i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_b_i_2_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_b_i_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_b_i_3_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_b_i_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_b_i_4_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_b_i_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_b_i_5_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_b_i_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_unsigned_a_0_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_unsigned_a_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_round_0_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_round_0_),
		.ccff_tail(cby_4__2__1_ccff_tail));

	cby_4__3_ cby_4__3_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_bottom_in(sb_4__2__0_chany_top_out[0:95]),
		.chany_top_in(sb_4__3__0_chany_bottom_out[0:95]),
		.ccff_head(sb_4__2__0_ccff_tail),
		.chany_bottom_out(cby_4__3__0_chany_bottom_out[0:95]),
		.chany_top_out(cby_4__3__0_chany_top_out[0:95]),
		.left_grid_right_width_0_height_1_subtile_0__pin_a_i_8_(cby_4__3__0_left_grid_right_width_0_height_1_subtile_0__pin_a_i_8_),
		.left_grid_right_width_0_height_1_subtile_0__pin_a_i_9_(cby_4__3__0_left_grid_right_width_0_height_1_subtile_0__pin_a_i_9_),
		.left_grid_right_width_0_height_1_subtile_0__pin_a_i_10_(cby_4__3__0_left_grid_right_width_0_height_1_subtile_0__pin_a_i_10_),
		.left_grid_right_width_0_height_1_subtile_0__pin_a_i_11_(cby_4__3__0_left_grid_right_width_0_height_1_subtile_0__pin_a_i_11_),
		.left_grid_right_width_0_height_1_subtile_0__pin_a_i_12_(cby_4__3__0_left_grid_right_width_0_height_1_subtile_0__pin_a_i_12_),
		.left_grid_right_width_0_height_1_subtile_0__pin_a_i_13_(cby_4__3__0_left_grid_right_width_0_height_1_subtile_0__pin_a_i_13_),
		.left_grid_right_width_0_height_1_subtile_0__pin_acc_fir_i_3_(cby_4__3__0_left_grid_right_width_0_height_1_subtile_0__pin_acc_fir_i_3_),
		.left_grid_right_width_0_height_1_subtile_0__pin_acc_fir_i_4_(cby_4__3__0_left_grid_right_width_0_height_1_subtile_0__pin_acc_fir_i_4_),
		.left_grid_right_width_0_height_1_subtile_0__pin_b_i_6_(cby_4__3__0_left_grid_right_width_0_height_1_subtile_0__pin_b_i_6_),
		.left_grid_right_width_0_height_1_subtile_0__pin_b_i_7_(cby_4__3__0_left_grid_right_width_0_height_1_subtile_0__pin_b_i_7_),
		.left_grid_right_width_0_height_1_subtile_0__pin_b_i_8_(cby_4__3__0_left_grid_right_width_0_height_1_subtile_0__pin_b_i_8_),
		.left_grid_right_width_0_height_1_subtile_0__pin_b_i_9_(cby_4__3__0_left_grid_right_width_0_height_1_subtile_0__pin_b_i_9_),
		.left_grid_right_width_0_height_1_subtile_0__pin_b_i_10_(cby_4__3__0_left_grid_right_width_0_height_1_subtile_0__pin_b_i_10_),
		.left_grid_right_width_0_height_1_subtile_0__pin_b_i_11_(cby_4__3__0_left_grid_right_width_0_height_1_subtile_0__pin_b_i_11_),
		.left_grid_right_width_0_height_1_subtile_0__pin_unsigned_b_0_(cby_4__3__0_left_grid_right_width_0_height_1_subtile_0__pin_unsigned_b_0_),
		.left_grid_right_width_0_height_1_subtile_0__pin_subtract_0_(cby_4__3__0_left_grid_right_width_0_height_1_subtile_0__pin_subtract_0_),
		.ccff_tail(cby_4__3__0_ccff_tail));

	cby_4__3_ cby_4__6_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_bottom_in(sb_4__2__1_chany_top_out[0:95]),
		.chany_top_in(sb_4__3__1_chany_bottom_out[0:95]),
		.ccff_head(sb_4__2__1_ccff_tail),
		.chany_bottom_out(cby_4__3__1_chany_bottom_out[0:95]),
		.chany_top_out(cby_4__3__1_chany_top_out[0:95]),
		.left_grid_right_width_0_height_1_subtile_0__pin_a_i_8_(cby_4__3__1_left_grid_right_width_0_height_1_subtile_0__pin_a_i_8_),
		.left_grid_right_width_0_height_1_subtile_0__pin_a_i_9_(cby_4__3__1_left_grid_right_width_0_height_1_subtile_0__pin_a_i_9_),
		.left_grid_right_width_0_height_1_subtile_0__pin_a_i_10_(cby_4__3__1_left_grid_right_width_0_height_1_subtile_0__pin_a_i_10_),
		.left_grid_right_width_0_height_1_subtile_0__pin_a_i_11_(cby_4__3__1_left_grid_right_width_0_height_1_subtile_0__pin_a_i_11_),
		.left_grid_right_width_0_height_1_subtile_0__pin_a_i_12_(cby_4__3__1_left_grid_right_width_0_height_1_subtile_0__pin_a_i_12_),
		.left_grid_right_width_0_height_1_subtile_0__pin_a_i_13_(cby_4__3__1_left_grid_right_width_0_height_1_subtile_0__pin_a_i_13_),
		.left_grid_right_width_0_height_1_subtile_0__pin_acc_fir_i_3_(cby_4__3__1_left_grid_right_width_0_height_1_subtile_0__pin_acc_fir_i_3_),
		.left_grid_right_width_0_height_1_subtile_0__pin_acc_fir_i_4_(cby_4__3__1_left_grid_right_width_0_height_1_subtile_0__pin_acc_fir_i_4_),
		.left_grid_right_width_0_height_1_subtile_0__pin_b_i_6_(cby_4__3__1_left_grid_right_width_0_height_1_subtile_0__pin_b_i_6_),
		.left_grid_right_width_0_height_1_subtile_0__pin_b_i_7_(cby_4__3__1_left_grid_right_width_0_height_1_subtile_0__pin_b_i_7_),
		.left_grid_right_width_0_height_1_subtile_0__pin_b_i_8_(cby_4__3__1_left_grid_right_width_0_height_1_subtile_0__pin_b_i_8_),
		.left_grid_right_width_0_height_1_subtile_0__pin_b_i_9_(cby_4__3__1_left_grid_right_width_0_height_1_subtile_0__pin_b_i_9_),
		.left_grid_right_width_0_height_1_subtile_0__pin_b_i_10_(cby_4__3__1_left_grid_right_width_0_height_1_subtile_0__pin_b_i_10_),
		.left_grid_right_width_0_height_1_subtile_0__pin_b_i_11_(cby_4__3__1_left_grid_right_width_0_height_1_subtile_0__pin_b_i_11_),
		.left_grid_right_width_0_height_1_subtile_0__pin_unsigned_b_0_(cby_4__3__1_left_grid_right_width_0_height_1_subtile_0__pin_unsigned_b_0_),
		.left_grid_right_width_0_height_1_subtile_0__pin_subtract_0_(cby_4__3__1_left_grid_right_width_0_height_1_subtile_0__pin_subtract_0_),
		.ccff_tail(cby_4__3__1_ccff_tail));

	cby_4__4_ cby_4__4_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_bottom_in(sb_4__3__0_chany_top_out[0:95]),
		.chany_top_in(sb_4__4__0_chany_bottom_out[0:95]),
		.ccff_head(sb_4__3__0_ccff_tail),
		.chany_bottom_out(cby_4__4__0_chany_bottom_out[0:95]),
		.chany_top_out(cby_4__4__0_chany_top_out[0:95]),
		.left_grid_right_width_0_height_2_subtile_0__pin_a_i_14_(cby_4__4__0_left_grid_right_width_0_height_2_subtile_0__pin_a_i_14_),
		.left_grid_right_width_0_height_2_subtile_0__pin_a_i_15_(cby_4__4__0_left_grid_right_width_0_height_2_subtile_0__pin_a_i_15_),
		.left_grid_right_width_0_height_2_subtile_0__pin_a_i_16_(cby_4__4__0_left_grid_right_width_0_height_2_subtile_0__pin_a_i_16_),
		.left_grid_right_width_0_height_2_subtile_0__pin_a_i_17_(cby_4__4__0_left_grid_right_width_0_height_2_subtile_0__pin_a_i_17_),
		.left_grid_right_width_0_height_2_subtile_0__pin_a_i_18_(cby_4__4__0_left_grid_right_width_0_height_2_subtile_0__pin_a_i_18_),
		.left_grid_right_width_0_height_2_subtile_0__pin_a_i_19_(cby_4__4__0_left_grid_right_width_0_height_2_subtile_0__pin_a_i_19_),
		.left_grid_right_width_0_height_2_subtile_0__pin_acc_fir_i_5_(cby_4__4__0_left_grid_right_width_0_height_2_subtile_0__pin_acc_fir_i_5_),
		.left_grid_right_width_0_height_2_subtile_0__pin_b_i_12_(cby_4__4__0_left_grid_right_width_0_height_2_subtile_0__pin_b_i_12_),
		.left_grid_right_width_0_height_2_subtile_0__pin_b_i_13_(cby_4__4__0_left_grid_right_width_0_height_2_subtile_0__pin_b_i_13_),
		.left_grid_right_width_0_height_2_subtile_0__pin_b_i_14_(cby_4__4__0_left_grid_right_width_0_height_2_subtile_0__pin_b_i_14_),
		.left_grid_right_width_0_height_2_subtile_0__pin_b_i_15_(cby_4__4__0_left_grid_right_width_0_height_2_subtile_0__pin_b_i_15_),
		.left_grid_right_width_0_height_2_subtile_0__pin_b_i_16_(cby_4__4__0_left_grid_right_width_0_height_2_subtile_0__pin_b_i_16_),
		.left_grid_right_width_0_height_2_subtile_0__pin_b_i_17_(cby_4__4__0_left_grid_right_width_0_height_2_subtile_0__pin_b_i_17_),
		.left_grid_right_width_0_height_2_subtile_0__pin_load_acc_0_(cby_4__4__0_left_grid_right_width_0_height_2_subtile_0__pin_load_acc_0_),
		.left_grid_right_width_0_height_2_subtile_0__pin_saturate_enable_0_(cby_4__4__0_left_grid_right_width_0_height_2_subtile_0__pin_saturate_enable_0_),
		.ccff_tail(cby_4__4__0_ccff_tail));

	cby_4__4_ cby_4__7_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_bottom_in(sb_4__3__1_chany_top_out[0:95]),
		.chany_top_in(sb_4__7__0_chany_bottom_out[0:95]),
		.ccff_head(sb_4__3__1_ccff_tail),
		.chany_bottom_out(cby_4__4__1_chany_bottom_out[0:95]),
		.chany_top_out(cby_4__4__1_chany_top_out[0:95]),
		.left_grid_right_width_0_height_2_subtile_0__pin_a_i_14_(cby_4__4__1_left_grid_right_width_0_height_2_subtile_0__pin_a_i_14_),
		.left_grid_right_width_0_height_2_subtile_0__pin_a_i_15_(cby_4__4__1_left_grid_right_width_0_height_2_subtile_0__pin_a_i_15_),
		.left_grid_right_width_0_height_2_subtile_0__pin_a_i_16_(cby_4__4__1_left_grid_right_width_0_height_2_subtile_0__pin_a_i_16_),
		.left_grid_right_width_0_height_2_subtile_0__pin_a_i_17_(cby_4__4__1_left_grid_right_width_0_height_2_subtile_0__pin_a_i_17_),
		.left_grid_right_width_0_height_2_subtile_0__pin_a_i_18_(cby_4__4__1_left_grid_right_width_0_height_2_subtile_0__pin_a_i_18_),
		.left_grid_right_width_0_height_2_subtile_0__pin_a_i_19_(cby_4__4__1_left_grid_right_width_0_height_2_subtile_0__pin_a_i_19_),
		.left_grid_right_width_0_height_2_subtile_0__pin_acc_fir_i_5_(cby_4__4__1_left_grid_right_width_0_height_2_subtile_0__pin_acc_fir_i_5_),
		.left_grid_right_width_0_height_2_subtile_0__pin_b_i_12_(cby_4__4__1_left_grid_right_width_0_height_2_subtile_0__pin_b_i_12_),
		.left_grid_right_width_0_height_2_subtile_0__pin_b_i_13_(cby_4__4__1_left_grid_right_width_0_height_2_subtile_0__pin_b_i_13_),
		.left_grid_right_width_0_height_2_subtile_0__pin_b_i_14_(cby_4__4__1_left_grid_right_width_0_height_2_subtile_0__pin_b_i_14_),
		.left_grid_right_width_0_height_2_subtile_0__pin_b_i_15_(cby_4__4__1_left_grid_right_width_0_height_2_subtile_0__pin_b_i_15_),
		.left_grid_right_width_0_height_2_subtile_0__pin_b_i_16_(cby_4__4__1_left_grid_right_width_0_height_2_subtile_0__pin_b_i_16_),
		.left_grid_right_width_0_height_2_subtile_0__pin_b_i_17_(cby_4__4__1_left_grid_right_width_0_height_2_subtile_0__pin_b_i_17_),
		.left_grid_right_width_0_height_2_subtile_0__pin_load_acc_0_(cby_4__4__1_left_grid_right_width_0_height_2_subtile_0__pin_load_acc_0_),
		.left_grid_right_width_0_height_2_subtile_0__pin_saturate_enable_0_(cby_4__4__1_left_grid_right_width_0_height_2_subtile_0__pin_saturate_enable_0_),
		.ccff_tail(cby_4__4__1_ccff_tail));

	cby_7__2_ cby_7__2_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_bottom_in(sb_7__1__0_chany_top_out[0:95]),
		.chany_top_in(sb_7__2__0_chany_bottom_out[0:95]),
		.ccff_head(cbx_7__1__0_ccff_tail),
		.chany_bottom_out(cby_7__2__0_chany_bottom_out[0:95]),
		.chany_top_out(cby_7__2__0_chany_top_out[0:95]),
		.left_grid_right_width_0_height_0_subtile_0__pin_ADDR_A1_i_2_(cby_7__2__0_left_grid_right_width_0_height_0_subtile_0__pin_ADDR_A1_i_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ADDR_A1_i_3_(cby_7__2__0_left_grid_right_width_0_height_0_subtile_0__pin_ADDR_A1_i_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ADDR_A1_i_4_(cby_7__2__0_left_grid_right_width_0_height_0_subtile_0__pin_ADDR_A1_i_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ADDR_A1_i_5_(cby_7__2__0_left_grid_right_width_0_height_0_subtile_0__pin_ADDR_A1_i_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_WDATA_B1_i_1_(cby_7__2__0_left_grid_right_width_0_height_0_subtile_0__pin_WDATA_B1_i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_WDATA_B1_i_2_(cby_7__2__0_left_grid_right_width_0_height_0_subtile_0__pin_WDATA_B1_i_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_WDATA_B1_i_3_(cby_7__2__0_left_grid_right_width_0_height_0_subtile_0__pin_WDATA_B1_i_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_WDATA_B1_i_4_(cby_7__2__0_left_grid_right_width_0_height_0_subtile_0__pin_WDATA_B1_i_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_WDATA_B1_i_5_(cby_7__2__0_left_grid_right_width_0_height_0_subtile_0__pin_WDATA_B1_i_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_WDATA_B1_i_6_(cby_7__2__0_left_grid_right_width_0_height_0_subtile_0__pin_WDATA_B1_i_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_WDATA_B1_i_7_(cby_7__2__0_left_grid_right_width_0_height_0_subtile_0__pin_WDATA_B1_i_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_WDATA_B1_i_8_(cby_7__2__0_left_grid_right_width_0_height_0_subtile_0__pin_WDATA_B1_i_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_WDATA_B1_i_9_(cby_7__2__0_left_grid_right_width_0_height_0_subtile_0__pin_WDATA_B1_i_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_WDATA_B1_i_10_(cby_7__2__0_left_grid_right_width_0_height_0_subtile_0__pin_WDATA_B1_i_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_WDATA_B1_i_11_(cby_7__2__0_left_grid_right_width_0_height_0_subtile_0__pin_WDATA_B1_i_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_WDATA_B1_i_12_(cby_7__2__0_left_grid_right_width_0_height_0_subtile_0__pin_WDATA_B1_i_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_WDATA_B1_i_13_(cby_7__2__0_left_grid_right_width_0_height_0_subtile_0__pin_WDATA_B1_i_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_WDATA_B1_i_14_(cby_7__2__0_left_grid_right_width_0_height_0_subtile_0__pin_WDATA_B1_i_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_WDATA_B1_i_15_(cby_7__2__0_left_grid_right_width_0_height_0_subtile_0__pin_WDATA_B1_i_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_WDATA_B1_i_16_(cby_7__2__0_left_grid_right_width_0_height_0_subtile_0__pin_WDATA_B1_i_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ADDR_B1_i_0_(cby_7__2__0_left_grid_right_width_0_height_0_subtile_0__pin_ADDR_B1_i_0_),
		.ccff_tail(cby_7__2__0_ccff_tail));

	cby_7__3_ cby_7__3_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_bottom_in(sb_7__2__0_chany_top_out[0:95]),
		.chany_top_in(sb_7__2__1_chany_bottom_out[0:95]),
		.ccff_head(sb_7__2__0_ccff_tail),
		.chany_bottom_out(cby_7__3__0_chany_bottom_out[0:95]),
		.chany_top_out(cby_7__3__0_chany_top_out[0:95]),
		.left_grid_right_width_0_height_1_subtile_0__pin_WDATA_A2_i_17_(cby_7__3__0_left_grid_right_width_0_height_1_subtile_0__pin_WDATA_A2_i_17_),
		.left_grid_right_width_0_height_1_subtile_0__pin_ADDR_A2_i_1_(cby_7__3__0_left_grid_right_width_0_height_1_subtile_0__pin_ADDR_A2_i_1_),
		.left_grid_right_width_0_height_1_subtile_0__pin_REN_A1_i_0_(cby_7__3__0_left_grid_right_width_0_height_1_subtile_0__pin_REN_A1_i_0_),
		.left_grid_right_width_0_height_1_subtile_0__pin_REN_A2_i_0_(cby_7__3__0_left_grid_right_width_0_height_1_subtile_0__pin_REN_A2_i_0_),
		.left_grid_right_width_0_height_1_subtile_0__pin_WEN_A2_i_0_(cby_7__3__0_left_grid_right_width_0_height_1_subtile_0__pin_WEN_A2_i_0_),
		.left_grid_right_width_0_height_1_subtile_0__pin_BE_A2_i_0_(cby_7__3__0_left_grid_right_width_0_height_1_subtile_0__pin_BE_A2_i_0_),
		.left_grid_right_width_0_height_1_subtile_0__pin_BE_A2_i_1_(cby_7__3__0_left_grid_right_width_0_height_1_subtile_0__pin_BE_A2_i_1_),
		.left_grid_right_width_0_height_1_subtile_0__pin_WDATA_B1_i_0_(cby_7__3__0_left_grid_right_width_0_height_1_subtile_0__pin_WDATA_B1_i_0_),
		.left_grid_right_width_0_height_1_subtile_0__pin_ADDR_B1_i_2_(cby_7__3__0_left_grid_right_width_0_height_1_subtile_0__pin_ADDR_B1_i_2_),
		.left_grid_right_width_0_height_1_subtile_0__pin_ADDR_B1_i_3_(cby_7__3__0_left_grid_right_width_0_height_1_subtile_0__pin_ADDR_B1_i_3_),
		.left_grid_right_width_0_height_1_subtile_0__pin_ADDR_B1_i_4_(cby_7__3__0_left_grid_right_width_0_height_1_subtile_0__pin_ADDR_B1_i_4_),
		.left_grid_right_width_0_height_1_subtile_0__pin_ADDR_B1_i_5_(cby_7__3__0_left_grid_right_width_0_height_1_subtile_0__pin_ADDR_B1_i_5_),
		.left_grid_right_width_0_height_1_subtile_0__pin_ADDR_B1_i_6_(cby_7__3__0_left_grid_right_width_0_height_1_subtile_0__pin_ADDR_B1_i_6_),
		.left_grid_right_width_0_height_1_subtile_0__pin_ADDR_B1_i_7_(cby_7__3__0_left_grid_right_width_0_height_1_subtile_0__pin_ADDR_B1_i_7_),
		.left_grid_right_width_0_height_1_subtile_0__pin_ADDR_B1_i_8_(cby_7__3__0_left_grid_right_width_0_height_1_subtile_0__pin_ADDR_B1_i_8_),
		.left_grid_right_width_0_height_1_subtile_0__pin_ADDR_B1_i_9_(cby_7__3__0_left_grid_right_width_0_height_1_subtile_0__pin_ADDR_B1_i_9_),
		.left_grid_right_width_0_height_1_subtile_0__pin_ADDR_B1_i_10_(cby_7__3__0_left_grid_right_width_0_height_1_subtile_0__pin_ADDR_B1_i_10_),
		.left_grid_right_width_0_height_1_subtile_0__pin_ADDR_B1_i_11_(cby_7__3__0_left_grid_right_width_0_height_1_subtile_0__pin_ADDR_B1_i_11_),
		.left_grid_right_width_0_height_1_subtile_0__pin_ADDR_B1_i_12_(cby_7__3__0_left_grid_right_width_0_height_1_subtile_0__pin_ADDR_B1_i_12_),
		.left_grid_right_width_0_height_1_subtile_0__pin_ADDR_B1_i_13_(cby_7__3__0_left_grid_right_width_0_height_1_subtile_0__pin_ADDR_B1_i_13_),
		.left_grid_right_width_0_height_1_subtile_0__pin_ADDR_B1_i_14_(cby_7__3__0_left_grid_right_width_0_height_1_subtile_0__pin_ADDR_B1_i_14_),
		.left_grid_right_width_0_height_1_subtile_0__pin_FLUSH2_i_0_(cby_7__3__0_left_grid_right_width_0_height_1_subtile_0__pin_FLUSH2_i_0_),
		.ccff_tail(cby_7__3__0_ccff_tail));

	cby_7__4_ cby_7__4_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_bottom_in(sb_7__2__1_chany_top_out[0:95]),
		.chany_top_in(sb_7__2__2_chany_bottom_out[0:95]),
		.ccff_head(sb_7__2__1_ccff_tail),
		.chany_bottom_out(cby_7__4__0_chany_bottom_out[0:95]),
		.chany_top_out(cby_7__4__0_chany_top_out[0:95]),
		.left_grid_right_width_0_height_2_subtile_0__pin_WDATA_A2_i_9_(cby_7__4__0_left_grid_right_width_0_height_2_subtile_0__pin_WDATA_A2_i_9_),
		.left_grid_right_width_0_height_2_subtile_0__pin_WDATA_A2_i_10_(cby_7__4__0_left_grid_right_width_0_height_2_subtile_0__pin_WDATA_A2_i_10_),
		.left_grid_right_width_0_height_2_subtile_0__pin_WDATA_A2_i_11_(cby_7__4__0_left_grid_right_width_0_height_2_subtile_0__pin_WDATA_A2_i_11_),
		.left_grid_right_width_0_height_2_subtile_0__pin_WDATA_A2_i_12_(cby_7__4__0_left_grid_right_width_0_height_2_subtile_0__pin_WDATA_A2_i_12_),
		.left_grid_right_width_0_height_2_subtile_0__pin_WDATA_A2_i_13_(cby_7__4__0_left_grid_right_width_0_height_2_subtile_0__pin_WDATA_A2_i_13_),
		.left_grid_right_width_0_height_2_subtile_0__pin_WDATA_A2_i_14_(cby_7__4__0_left_grid_right_width_0_height_2_subtile_0__pin_WDATA_A2_i_14_),
		.left_grid_right_width_0_height_2_subtile_0__pin_WDATA_A2_i_15_(cby_7__4__0_left_grid_right_width_0_height_2_subtile_0__pin_WDATA_A2_i_15_),
		.left_grid_right_width_0_height_2_subtile_0__pin_WDATA_A2_i_16_(cby_7__4__0_left_grid_right_width_0_height_2_subtile_0__pin_WDATA_A2_i_16_),
		.left_grid_right_width_0_height_2_subtile_0__pin_ADDR_A2_i_0_(cby_7__4__0_left_grid_right_width_0_height_2_subtile_0__pin_ADDR_A2_i_0_),
		.left_grid_right_width_0_height_2_subtile_0__pin_ADDR_A2_i_2_(cby_7__4__0_left_grid_right_width_0_height_2_subtile_0__pin_ADDR_A2_i_2_),
		.left_grid_right_width_0_height_2_subtile_0__pin_ADDR_A2_i_3_(cby_7__4__0_left_grid_right_width_0_height_2_subtile_0__pin_ADDR_A2_i_3_),
		.left_grid_right_width_0_height_2_subtile_0__pin_ADDR_A2_i_4_(cby_7__4__0_left_grid_right_width_0_height_2_subtile_0__pin_ADDR_A2_i_4_),
		.left_grid_right_width_0_height_2_subtile_0__pin_ADDR_A2_i_5_(cby_7__4__0_left_grid_right_width_0_height_2_subtile_0__pin_ADDR_A2_i_5_),
		.left_grid_right_width_0_height_2_subtile_0__pin_ADDR_A2_i_6_(cby_7__4__0_left_grid_right_width_0_height_2_subtile_0__pin_ADDR_A2_i_6_),
		.left_grid_right_width_0_height_2_subtile_0__pin_ADDR_A2_i_7_(cby_7__4__0_left_grid_right_width_0_height_2_subtile_0__pin_ADDR_A2_i_7_),
		.left_grid_right_width_0_height_2_subtile_0__pin_ADDR_A2_i_8_(cby_7__4__0_left_grid_right_width_0_height_2_subtile_0__pin_ADDR_A2_i_8_),
		.left_grid_right_width_0_height_2_subtile_0__pin_ADDR_A2_i_9_(cby_7__4__0_left_grid_right_width_0_height_2_subtile_0__pin_ADDR_A2_i_9_),
		.left_grid_right_width_0_height_2_subtile_0__pin_ADDR_A2_i_10_(cby_7__4__0_left_grid_right_width_0_height_2_subtile_0__pin_ADDR_A2_i_10_),
		.left_grid_right_width_0_height_2_subtile_0__pin_ADDR_A2_i_11_(cby_7__4__0_left_grid_right_width_0_height_2_subtile_0__pin_ADDR_A2_i_11_),
		.left_grid_right_width_0_height_2_subtile_0__pin_ADDR_A2_i_12_(cby_7__4__0_left_grid_right_width_0_height_2_subtile_0__pin_ADDR_A2_i_12_),
		.left_grid_right_width_0_height_2_subtile_0__pin_ADDR_A2_i_13_(cby_7__4__0_left_grid_right_width_0_height_2_subtile_0__pin_ADDR_A2_i_13_),
		.left_grid_right_width_0_height_2_subtile_0__pin_WEN_A1_i_0_(cby_7__4__0_left_grid_right_width_0_height_2_subtile_0__pin_WEN_A1_i_0_),
		.ccff_tail(cby_7__4__0_ccff_tail));

	cby_7__5_ cby_7__5_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_bottom_in(sb_7__2__2_chany_top_out[0:95]),
		.chany_top_in(sb_7__2__3_chany_bottom_out[0:95]),
		.ccff_head(sb_7__2__2_ccff_tail),
		.chany_bottom_out(cby_7__5__0_chany_bottom_out[0:95]),
		.chany_top_out(cby_7__5__0_chany_top_out[0:95]),
		.left_grid_right_width_0_height_3_subtile_0__pin_WDATA_A1_i_7_(cby_7__5__0_left_grid_right_width_0_height_3_subtile_0__pin_WDATA_A1_i_7_),
		.left_grid_right_width_0_height_3_subtile_0__pin_WDATA_A1_i_8_(cby_7__5__0_left_grid_right_width_0_height_3_subtile_0__pin_WDATA_A1_i_8_),
		.left_grid_right_width_0_height_3_subtile_0__pin_WDATA_A1_i_9_(cby_7__5__0_left_grid_right_width_0_height_3_subtile_0__pin_WDATA_A1_i_9_),
		.left_grid_right_width_0_height_3_subtile_0__pin_WDATA_A1_i_10_(cby_7__5__0_left_grid_right_width_0_height_3_subtile_0__pin_WDATA_A1_i_10_),
		.left_grid_right_width_0_height_3_subtile_0__pin_WDATA_A1_i_11_(cby_7__5__0_left_grid_right_width_0_height_3_subtile_0__pin_WDATA_A1_i_11_),
		.left_grid_right_width_0_height_3_subtile_0__pin_WDATA_A1_i_12_(cby_7__5__0_left_grid_right_width_0_height_3_subtile_0__pin_WDATA_A1_i_12_),
		.left_grid_right_width_0_height_3_subtile_0__pin_WDATA_A1_i_13_(cby_7__5__0_left_grid_right_width_0_height_3_subtile_0__pin_WDATA_A1_i_13_),
		.left_grid_right_width_0_height_3_subtile_0__pin_WDATA_A1_i_14_(cby_7__5__0_left_grid_right_width_0_height_3_subtile_0__pin_WDATA_A1_i_14_),
		.left_grid_right_width_0_height_3_subtile_0__pin_WDATA_A1_i_15_(cby_7__5__0_left_grid_right_width_0_height_3_subtile_0__pin_WDATA_A1_i_15_),
		.left_grid_right_width_0_height_3_subtile_0__pin_WDATA_A1_i_16_(cby_7__5__0_left_grid_right_width_0_height_3_subtile_0__pin_WDATA_A1_i_16_),
		.left_grid_right_width_0_height_3_subtile_0__pin_WDATA_A1_i_17_(cby_7__5__0_left_grid_right_width_0_height_3_subtile_0__pin_WDATA_A1_i_17_),
		.left_grid_right_width_0_height_3_subtile_0__pin_ADDR_A1_i_0_(cby_7__5__0_left_grid_right_width_0_height_3_subtile_0__pin_ADDR_A1_i_0_),
		.left_grid_right_width_0_height_3_subtile_0__pin_ADDR_A1_i_1_(cby_7__5__0_left_grid_right_width_0_height_3_subtile_0__pin_ADDR_A1_i_1_),
		.left_grid_right_width_0_height_3_subtile_0__pin_BE_A1_i_0_(cby_7__5__0_left_grid_right_width_0_height_3_subtile_0__pin_BE_A1_i_0_),
		.left_grid_right_width_0_height_3_subtile_0__pin_BE_A1_i_1_(cby_7__5__0_left_grid_right_width_0_height_3_subtile_0__pin_BE_A1_i_1_),
		.left_grid_right_width_0_height_3_subtile_0__pin_REN_B2_i_0_(cby_7__5__0_left_grid_right_width_0_height_3_subtile_0__pin_REN_B2_i_0_),
		.left_grid_right_width_0_height_3_subtile_0__pin_WEN_B2_i_0_(cby_7__5__0_left_grid_right_width_0_height_3_subtile_0__pin_WEN_B2_i_0_),
		.left_grid_right_width_0_height_3_subtile_0__pin_BE_B1_i_0_(cby_7__5__0_left_grid_right_width_0_height_3_subtile_0__pin_BE_B1_i_0_),
		.left_grid_right_width_0_height_3_subtile_0__pin_BE_B1_i_1_(cby_7__5__0_left_grid_right_width_0_height_3_subtile_0__pin_BE_B1_i_1_),
		.left_grid_right_width_0_height_3_subtile_0__pin_BE_B2_i_0_(cby_7__5__0_left_grid_right_width_0_height_3_subtile_0__pin_BE_B2_i_0_),
		.left_grid_right_width_0_height_3_subtile_0__pin_BE_B2_i_1_(cby_7__5__0_left_grid_right_width_0_height_3_subtile_0__pin_BE_B2_i_1_),
		.left_grid_right_width_0_height_3_subtile_0__pin_FLUSH1_i_0_(cby_7__5__0_left_grid_right_width_0_height_3_subtile_0__pin_FLUSH1_i_0_),
		.ccff_tail(cby_7__5__0_ccff_tail));

	cby_7__6_ cby_7__6_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_bottom_in(sb_7__2__3_chany_top_out[0:95]),
		.chany_top_in(sb_7__2__4_chany_bottom_out[0:95]),
		.ccff_head(sb_7__2__3_ccff_tail),
		.chany_bottom_out(cby_7__6__0_chany_bottom_out[0:95]),
		.chany_top_out(cby_7__6__0_chany_top_out[0:95]),
		.left_grid_right_width_0_height_4_subtile_0__pin_WDATA_A2_i_0_(cby_7__6__0_left_grid_right_width_0_height_4_subtile_0__pin_WDATA_A2_i_0_),
		.left_grid_right_width_0_height_4_subtile_0__pin_WDATA_A2_i_1_(cby_7__6__0_left_grid_right_width_0_height_4_subtile_0__pin_WDATA_A2_i_1_),
		.left_grid_right_width_0_height_4_subtile_0__pin_WDATA_A2_i_2_(cby_7__6__0_left_grid_right_width_0_height_4_subtile_0__pin_WDATA_A2_i_2_),
		.left_grid_right_width_0_height_4_subtile_0__pin_WDATA_A2_i_3_(cby_7__6__0_left_grid_right_width_0_height_4_subtile_0__pin_WDATA_A2_i_3_),
		.left_grid_right_width_0_height_4_subtile_0__pin_WDATA_A2_i_4_(cby_7__6__0_left_grid_right_width_0_height_4_subtile_0__pin_WDATA_A2_i_4_),
		.left_grid_right_width_0_height_4_subtile_0__pin_WDATA_A2_i_5_(cby_7__6__0_left_grid_right_width_0_height_4_subtile_0__pin_WDATA_A2_i_5_),
		.left_grid_right_width_0_height_4_subtile_0__pin_WDATA_A2_i_6_(cby_7__6__0_left_grid_right_width_0_height_4_subtile_0__pin_WDATA_A2_i_6_),
		.left_grid_right_width_0_height_4_subtile_0__pin_WDATA_A2_i_7_(cby_7__6__0_left_grid_right_width_0_height_4_subtile_0__pin_WDATA_A2_i_7_),
		.left_grid_right_width_0_height_4_subtile_0__pin_WDATA_A2_i_8_(cby_7__6__0_left_grid_right_width_0_height_4_subtile_0__pin_WDATA_A2_i_8_),
		.left_grid_right_width_0_height_4_subtile_0__pin_WDATA_B2_i_17_(cby_7__6__0_left_grid_right_width_0_height_4_subtile_0__pin_WDATA_B2_i_17_),
		.left_grid_right_width_0_height_4_subtile_0__pin_ADDR_B2_i_1_(cby_7__6__0_left_grid_right_width_0_height_4_subtile_0__pin_ADDR_B2_i_1_),
		.left_grid_right_width_0_height_4_subtile_0__pin_ADDR_B2_i_4_(cby_7__6__0_left_grid_right_width_0_height_4_subtile_0__pin_ADDR_B2_i_4_),
		.left_grid_right_width_0_height_4_subtile_0__pin_ADDR_B2_i_5_(cby_7__6__0_left_grid_right_width_0_height_4_subtile_0__pin_ADDR_B2_i_5_),
		.left_grid_right_width_0_height_4_subtile_0__pin_ADDR_B2_i_6_(cby_7__6__0_left_grid_right_width_0_height_4_subtile_0__pin_ADDR_B2_i_6_),
		.left_grid_right_width_0_height_4_subtile_0__pin_ADDR_B2_i_7_(cby_7__6__0_left_grid_right_width_0_height_4_subtile_0__pin_ADDR_B2_i_7_),
		.left_grid_right_width_0_height_4_subtile_0__pin_ADDR_B2_i_8_(cby_7__6__0_left_grid_right_width_0_height_4_subtile_0__pin_ADDR_B2_i_8_),
		.left_grid_right_width_0_height_4_subtile_0__pin_ADDR_B2_i_9_(cby_7__6__0_left_grid_right_width_0_height_4_subtile_0__pin_ADDR_B2_i_9_),
		.left_grid_right_width_0_height_4_subtile_0__pin_ADDR_B2_i_10_(cby_7__6__0_left_grid_right_width_0_height_4_subtile_0__pin_ADDR_B2_i_10_),
		.left_grid_right_width_0_height_4_subtile_0__pin_ADDR_B2_i_11_(cby_7__6__0_left_grid_right_width_0_height_4_subtile_0__pin_ADDR_B2_i_11_),
		.left_grid_right_width_0_height_4_subtile_0__pin_ADDR_B2_i_12_(cby_7__6__0_left_grid_right_width_0_height_4_subtile_0__pin_ADDR_B2_i_12_),
		.left_grid_right_width_0_height_4_subtile_0__pin_ADDR_B2_i_13_(cby_7__6__0_left_grid_right_width_0_height_4_subtile_0__pin_ADDR_B2_i_13_),
		.left_grid_right_width_0_height_4_subtile_0__pin_WEN_B1_i_0_(cby_7__6__0_left_grid_right_width_0_height_4_subtile_0__pin_WEN_B1_i_0_),
		.ccff_tail(cby_7__6__0_ccff_tail));

	cby_7__7_ cby_7__7_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_bottom_in(sb_7__2__4_chany_top_out[0:95]),
		.chany_top_in(sb_7__7__0_chany_bottom_out[0:95]),
		.ccff_head(sb_7__2__4_ccff_tail),
		.chany_bottom_out(cby_7__7__0_chany_bottom_out[0:95]),
		.chany_top_out(cby_7__7__0_chany_top_out[0:95]),
		.left_grid_right_width_0_height_5_subtile_0__pin_WDATA_B2_i_0_(cby_7__7__0_left_grid_right_width_0_height_5_subtile_0__pin_WDATA_B2_i_0_),
		.left_grid_right_width_0_height_5_subtile_0__pin_WDATA_B2_i_1_(cby_7__7__0_left_grid_right_width_0_height_5_subtile_0__pin_WDATA_B2_i_1_),
		.left_grid_right_width_0_height_5_subtile_0__pin_WDATA_B2_i_2_(cby_7__7__0_left_grid_right_width_0_height_5_subtile_0__pin_WDATA_B2_i_2_),
		.left_grid_right_width_0_height_5_subtile_0__pin_WDATA_B2_i_3_(cby_7__7__0_left_grid_right_width_0_height_5_subtile_0__pin_WDATA_B2_i_3_),
		.left_grid_right_width_0_height_5_subtile_0__pin_WDATA_B2_i_4_(cby_7__7__0_left_grid_right_width_0_height_5_subtile_0__pin_WDATA_B2_i_4_),
		.left_grid_right_width_0_height_5_subtile_0__pin_WDATA_B2_i_5_(cby_7__7__0_left_grid_right_width_0_height_5_subtile_0__pin_WDATA_B2_i_5_),
		.left_grid_right_width_0_height_5_subtile_0__pin_WDATA_B2_i_6_(cby_7__7__0_left_grid_right_width_0_height_5_subtile_0__pin_WDATA_B2_i_6_),
		.left_grid_right_width_0_height_5_subtile_0__pin_WDATA_B2_i_7_(cby_7__7__0_left_grid_right_width_0_height_5_subtile_0__pin_WDATA_B2_i_7_),
		.left_grid_right_width_0_height_5_subtile_0__pin_WDATA_B2_i_8_(cby_7__7__0_left_grid_right_width_0_height_5_subtile_0__pin_WDATA_B2_i_8_),
		.left_grid_right_width_0_height_5_subtile_0__pin_WDATA_B2_i_9_(cby_7__7__0_left_grid_right_width_0_height_5_subtile_0__pin_WDATA_B2_i_9_),
		.left_grid_right_width_0_height_5_subtile_0__pin_WDATA_B2_i_10_(cby_7__7__0_left_grid_right_width_0_height_5_subtile_0__pin_WDATA_B2_i_10_),
		.left_grid_right_width_0_height_5_subtile_0__pin_WDATA_B2_i_11_(cby_7__7__0_left_grid_right_width_0_height_5_subtile_0__pin_WDATA_B2_i_11_),
		.left_grid_right_width_0_height_5_subtile_0__pin_WDATA_B2_i_12_(cby_7__7__0_left_grid_right_width_0_height_5_subtile_0__pin_WDATA_B2_i_12_),
		.left_grid_right_width_0_height_5_subtile_0__pin_WDATA_B2_i_13_(cby_7__7__0_left_grid_right_width_0_height_5_subtile_0__pin_WDATA_B2_i_13_),
		.left_grid_right_width_0_height_5_subtile_0__pin_WDATA_B2_i_14_(cby_7__7__0_left_grid_right_width_0_height_5_subtile_0__pin_WDATA_B2_i_14_),
		.left_grid_right_width_0_height_5_subtile_0__pin_WDATA_B2_i_15_(cby_7__7__0_left_grid_right_width_0_height_5_subtile_0__pin_WDATA_B2_i_15_),
		.left_grid_right_width_0_height_5_subtile_0__pin_WDATA_B2_i_16_(cby_7__7__0_left_grid_right_width_0_height_5_subtile_0__pin_WDATA_B2_i_16_),
		.left_grid_right_width_0_height_5_subtile_0__pin_ADDR_B2_i_0_(cby_7__7__0_left_grid_right_width_0_height_5_subtile_0__pin_ADDR_B2_i_0_),
		.left_grid_right_width_0_height_5_subtile_0__pin_ADDR_B2_i_2_(cby_7__7__0_left_grid_right_width_0_height_5_subtile_0__pin_ADDR_B2_i_2_),
		.left_grid_right_width_0_height_5_subtile_0__pin_ADDR_B2_i_3_(cby_7__7__0_left_grid_right_width_0_height_5_subtile_0__pin_ADDR_B2_i_3_),
		.left_grid_right_width_0_height_5_subtile_0__pin_REN_B1_i_0_(cby_7__7__0_left_grid_right_width_0_height_5_subtile_0__pin_REN_B1_i_0_),
		.ccff_tail(cby_7__7__0_ccff_tail));

	cby_9__1_ cby_9__1_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_bottom_in(sb_1__0__1_chany_top_out[0:95]),
		.chany_top_in(sb_9__1__0_chany_bottom_out[0:95]),
		.ccff_head(sb_1__0__1_ccff_tail),
		.chany_bottom_out(cby_9__1__0_chany_bottom_out[0:95]),
		.chany_top_out(cby_9__1__0_chany_top_out[0:95]),
		.right_grid_left_width_0_height_0_subtile_0__pin_f2a_i_0_(cby_9__1__0_right_grid_left_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_f2a_i_0_(cby_9__1__0_right_grid_left_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_f2a_i_0_(cby_9__1__0_right_grid_left_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_f2a_i_0_(cby_9__1__0_right_grid_left_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_f2a_i_0_(cby_9__1__0_right_grid_left_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_f2a_i_0_(cby_9__1__0_right_grid_left_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_f2a_i_0_(cby_9__1__0_right_grid_left_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_f2a_i_0_(cby_9__1__0_right_grid_left_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_8__pin_f2a_i_0_(cby_9__1__0_right_grid_left_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_9__pin_f2a_i_0_(cby_9__1__0_right_grid_left_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_10__pin_f2a_i_0_(cby_9__1__0_right_grid_left_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_11__pin_f2a_i_0_(cby_9__1__0_right_grid_left_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_12__pin_f2a_i_0_(cby_9__1__0_right_grid_left_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_13__pin_f2a_i_0_(cby_9__1__0_right_grid_left_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_14__pin_f2a_i_0_(cby_9__1__0_right_grid_left_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_15__pin_f2a_i_0_(cby_9__1__0_right_grid_left_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_16__pin_f2a_i_0_(cby_9__1__0_right_grid_left_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_17__pin_f2a_i_0_(cby_9__1__0_right_grid_left_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_18__pin_f2a_i_0_(cby_9__1__0_right_grid_left_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_19__pin_f2a_i_0_(cby_9__1__0_right_grid_left_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.ccff_tail(cby_9__1__0_ccff_tail));

	cby_9__1_ cby_9__8_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_bottom_in(sb_9__7__0_chany_top_out[0:95]),
		.chany_top_in(sb_1__8__1_chany_bottom_out[0:95]),
		.ccff_head(cbx_2__7__5_ccff_tail),
		.chany_bottom_out(cby_9__1__1_chany_bottom_out[0:95]),
		.chany_top_out(cby_9__1__1_chany_top_out[0:95]),
		.right_grid_left_width_0_height_0_subtile_0__pin_f2a_i_0_(cby_9__1__1_right_grid_left_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_f2a_i_0_(cby_9__1__1_right_grid_left_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_f2a_i_0_(cby_9__1__1_right_grid_left_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_f2a_i_0_(cby_9__1__1_right_grid_left_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_f2a_i_0_(cby_9__1__1_right_grid_left_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_f2a_i_0_(cby_9__1__1_right_grid_left_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_f2a_i_0_(cby_9__1__1_right_grid_left_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_f2a_i_0_(cby_9__1__1_right_grid_left_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_8__pin_f2a_i_0_(cby_9__1__1_right_grid_left_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_9__pin_f2a_i_0_(cby_9__1__1_right_grid_left_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_10__pin_f2a_i_0_(cby_9__1__1_right_grid_left_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_11__pin_f2a_i_0_(cby_9__1__1_right_grid_left_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_12__pin_f2a_i_0_(cby_9__1__1_right_grid_left_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_13__pin_f2a_i_0_(cby_9__1__1_right_grid_left_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_14__pin_f2a_i_0_(cby_9__1__1_right_grid_left_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_15__pin_f2a_i_0_(cby_9__1__1_right_grid_left_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_16__pin_f2a_i_0_(cby_9__1__1_right_grid_left_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_17__pin_f2a_i_0_(cby_9__1__1_right_grid_left_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_18__pin_f2a_i_0_(cby_9__1__1_right_grid_left_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_19__pin_f2a_i_0_(cby_9__1__1_right_grid_left_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.ccff_tail(cby_9__1__1_ccff_tail));

	cby_9__2_ cby_9__2_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_bottom_in(sb_9__1__0_chany_top_out[0:95]),
		.chany_top_in(sb_9__2__0_chany_bottom_out[0:95]),
		.ccff_head(cbx_2__1__5_ccff_tail),
		.chany_bottom_out(cby_9__2__0_chany_bottom_out[0:95]),
		.chany_top_out(cby_9__2__0_chany_top_out[0:95]),
		.right_grid_left_width_0_height_0_subtile_0__pin_f2a_i_0_(cby_9__2__0_right_grid_left_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_f2a_i_0_(cby_9__2__0_right_grid_left_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_f2a_i_0_(cby_9__2__0_right_grid_left_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_f2a_i_0_(cby_9__2__0_right_grid_left_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_f2a_i_0_(cby_9__2__0_right_grid_left_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_f2a_i_0_(cby_9__2__0_right_grid_left_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_f2a_i_0_(cby_9__2__0_right_grid_left_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_f2a_i_0_(cby_9__2__0_right_grid_left_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_8__pin_f2a_i_0_(cby_9__2__0_right_grid_left_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_9__pin_f2a_i_0_(cby_9__2__0_right_grid_left_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_10__pin_f2a_i_0_(cby_9__2__0_right_grid_left_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_11__pin_f2a_i_0_(cby_9__2__0_right_grid_left_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_12__pin_f2a_i_0_(cby_9__2__0_right_grid_left_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_13__pin_f2a_i_0_(cby_9__2__0_right_grid_left_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_14__pin_f2a_i_0_(cby_9__2__0_right_grid_left_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_15__pin_f2a_i_0_(cby_9__2__0_right_grid_left_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_16__pin_f2a_i_0_(cby_9__2__0_right_grid_left_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_17__pin_f2a_i_0_(cby_9__2__0_right_grid_left_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_18__pin_f2a_i_0_(cby_9__2__0_right_grid_left_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_19__pin_f2a_i_0_(cby_9__2__0_right_grid_left_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_0_(cby_9__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_1_(cby_9__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_2_(cby_9__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_3_(cby_9__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_4_(cby_9__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_5_(cby_9__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_6_(cby_9__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_7_(cby_9__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_8_(cby_9__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_9_(cby_9__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_0_(cby_9__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_1_(cby_9__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_2_(cby_9__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_3_(cby_9__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_4_(cby_9__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_5_(cby_9__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_6_(cby_9__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_7_(cby_9__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_8_(cby_9__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_9_(cby_9__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_0_(cby_9__2__0_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_1_(cby_9__2__0_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_2_(cby_9__2__0_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_3_(cby_9__2__0_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_4_(cby_9__2__0_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_5_(cby_9__2__0_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.ccff_tail(cby_9__2__0_ccff_tail));

	cby_9__2_ cby_9__3_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_bottom_in(sb_9__2__0_chany_top_out[0:95]),
		.chany_top_in(sb_9__2__1_chany_bottom_out[0:95]),
		.ccff_head(cbx_2__2__25_ccff_tail),
		.chany_bottom_out(cby_9__2__1_chany_bottom_out[0:95]),
		.chany_top_out(cby_9__2__1_chany_top_out[0:95]),
		.right_grid_left_width_0_height_0_subtile_0__pin_f2a_i_0_(cby_9__2__1_right_grid_left_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_f2a_i_0_(cby_9__2__1_right_grid_left_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_f2a_i_0_(cby_9__2__1_right_grid_left_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_f2a_i_0_(cby_9__2__1_right_grid_left_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_f2a_i_0_(cby_9__2__1_right_grid_left_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_f2a_i_0_(cby_9__2__1_right_grid_left_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_f2a_i_0_(cby_9__2__1_right_grid_left_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_f2a_i_0_(cby_9__2__1_right_grid_left_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_8__pin_f2a_i_0_(cby_9__2__1_right_grid_left_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_9__pin_f2a_i_0_(cby_9__2__1_right_grid_left_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_10__pin_f2a_i_0_(cby_9__2__1_right_grid_left_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_11__pin_f2a_i_0_(cby_9__2__1_right_grid_left_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_12__pin_f2a_i_0_(cby_9__2__1_right_grid_left_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_13__pin_f2a_i_0_(cby_9__2__1_right_grid_left_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_14__pin_f2a_i_0_(cby_9__2__1_right_grid_left_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_15__pin_f2a_i_0_(cby_9__2__1_right_grid_left_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_16__pin_f2a_i_0_(cby_9__2__1_right_grid_left_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_17__pin_f2a_i_0_(cby_9__2__1_right_grid_left_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_18__pin_f2a_i_0_(cby_9__2__1_right_grid_left_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_19__pin_f2a_i_0_(cby_9__2__1_right_grid_left_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_0_(cby_9__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_1_(cby_9__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_2_(cby_9__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_3_(cby_9__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_4_(cby_9__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_5_(cby_9__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_6_(cby_9__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_7_(cby_9__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_8_(cby_9__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_9_(cby_9__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_0_(cby_9__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_1_(cby_9__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_2_(cby_9__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_3_(cby_9__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_4_(cby_9__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_5_(cby_9__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_6_(cby_9__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_7_(cby_9__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_8_(cby_9__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_9_(cby_9__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_0_(cby_9__2__1_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_1_(cby_9__2__1_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_2_(cby_9__2__1_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_3_(cby_9__2__1_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_4_(cby_9__2__1_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_5_(cby_9__2__1_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.ccff_tail(cby_9__2__1_ccff_tail));

	cby_9__2_ cby_9__4_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_bottom_in(sb_9__2__1_chany_top_out[0:95]),
		.chany_top_in(sb_9__2__2_chany_bottom_out[0:95]),
		.ccff_head(cbx_2__2__26_ccff_tail),
		.chany_bottom_out(cby_9__2__2_chany_bottom_out[0:95]),
		.chany_top_out(cby_9__2__2_chany_top_out[0:95]),
		.right_grid_left_width_0_height_0_subtile_0__pin_f2a_i_0_(cby_9__2__2_right_grid_left_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_f2a_i_0_(cby_9__2__2_right_grid_left_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_f2a_i_0_(cby_9__2__2_right_grid_left_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_f2a_i_0_(cby_9__2__2_right_grid_left_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_f2a_i_0_(cby_9__2__2_right_grid_left_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_f2a_i_0_(cby_9__2__2_right_grid_left_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_f2a_i_0_(cby_9__2__2_right_grid_left_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_f2a_i_0_(cby_9__2__2_right_grid_left_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_8__pin_f2a_i_0_(cby_9__2__2_right_grid_left_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_9__pin_f2a_i_0_(cby_9__2__2_right_grid_left_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_10__pin_f2a_i_0_(cby_9__2__2_right_grid_left_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_11__pin_f2a_i_0_(cby_9__2__2_right_grid_left_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_12__pin_f2a_i_0_(cby_9__2__2_right_grid_left_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_13__pin_f2a_i_0_(cby_9__2__2_right_grid_left_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_14__pin_f2a_i_0_(cby_9__2__2_right_grid_left_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_15__pin_f2a_i_0_(cby_9__2__2_right_grid_left_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_16__pin_f2a_i_0_(cby_9__2__2_right_grid_left_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_17__pin_f2a_i_0_(cby_9__2__2_right_grid_left_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_18__pin_f2a_i_0_(cby_9__2__2_right_grid_left_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_19__pin_f2a_i_0_(cby_9__2__2_right_grid_left_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_0_(cby_9__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_1_(cby_9__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_2_(cby_9__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_3_(cby_9__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_4_(cby_9__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_5_(cby_9__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_6_(cby_9__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_7_(cby_9__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_8_(cby_9__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_9_(cby_9__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_0_(cby_9__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_1_(cby_9__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_2_(cby_9__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_3_(cby_9__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_4_(cby_9__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_5_(cby_9__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_6_(cby_9__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_7_(cby_9__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_8_(cby_9__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_9_(cby_9__2__2_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_0_(cby_9__2__2_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_1_(cby_9__2__2_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_2_(cby_9__2__2_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_3_(cby_9__2__2_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_4_(cby_9__2__2_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_5_(cby_9__2__2_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.ccff_tail(cby_9__2__2_ccff_tail));

	cby_9__2_ cby_9__5_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_bottom_in(sb_9__2__2_chany_top_out[0:95]),
		.chany_top_in(sb_9__2__3_chany_bottom_out[0:95]),
		.ccff_head(cbx_2__2__27_ccff_tail),
		.chany_bottom_out(cby_9__2__3_chany_bottom_out[0:95]),
		.chany_top_out(cby_9__2__3_chany_top_out[0:95]),
		.right_grid_left_width_0_height_0_subtile_0__pin_f2a_i_0_(cby_9__2__3_right_grid_left_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_f2a_i_0_(cby_9__2__3_right_grid_left_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_f2a_i_0_(cby_9__2__3_right_grid_left_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_f2a_i_0_(cby_9__2__3_right_grid_left_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_f2a_i_0_(cby_9__2__3_right_grid_left_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_f2a_i_0_(cby_9__2__3_right_grid_left_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_f2a_i_0_(cby_9__2__3_right_grid_left_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_f2a_i_0_(cby_9__2__3_right_grid_left_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_8__pin_f2a_i_0_(cby_9__2__3_right_grid_left_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_9__pin_f2a_i_0_(cby_9__2__3_right_grid_left_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_10__pin_f2a_i_0_(cby_9__2__3_right_grid_left_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_11__pin_f2a_i_0_(cby_9__2__3_right_grid_left_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_12__pin_f2a_i_0_(cby_9__2__3_right_grid_left_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_13__pin_f2a_i_0_(cby_9__2__3_right_grid_left_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_14__pin_f2a_i_0_(cby_9__2__3_right_grid_left_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_15__pin_f2a_i_0_(cby_9__2__3_right_grid_left_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_16__pin_f2a_i_0_(cby_9__2__3_right_grid_left_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_17__pin_f2a_i_0_(cby_9__2__3_right_grid_left_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_18__pin_f2a_i_0_(cby_9__2__3_right_grid_left_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_19__pin_f2a_i_0_(cby_9__2__3_right_grid_left_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_0_(cby_9__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_1_(cby_9__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_2_(cby_9__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_3_(cby_9__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_4_(cby_9__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_5_(cby_9__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_6_(cby_9__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_7_(cby_9__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_8_(cby_9__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_9_(cby_9__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_0_(cby_9__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_1_(cby_9__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_2_(cby_9__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_3_(cby_9__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_4_(cby_9__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_5_(cby_9__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_6_(cby_9__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_7_(cby_9__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_8_(cby_9__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_9_(cby_9__2__3_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_0_(cby_9__2__3_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_1_(cby_9__2__3_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_2_(cby_9__2__3_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_3_(cby_9__2__3_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_4_(cby_9__2__3_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_5_(cby_9__2__3_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.ccff_tail(cby_9__2__3_ccff_tail));

	cby_9__2_ cby_9__6_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_bottom_in(sb_9__2__3_chany_top_out[0:95]),
		.chany_top_in(sb_9__2__4_chany_bottom_out[0:95]),
		.ccff_head(cbx_2__2__28_ccff_tail),
		.chany_bottom_out(cby_9__2__4_chany_bottom_out[0:95]),
		.chany_top_out(cby_9__2__4_chany_top_out[0:95]),
		.right_grid_left_width_0_height_0_subtile_0__pin_f2a_i_0_(cby_9__2__4_right_grid_left_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_f2a_i_0_(cby_9__2__4_right_grid_left_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_f2a_i_0_(cby_9__2__4_right_grid_left_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_f2a_i_0_(cby_9__2__4_right_grid_left_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_f2a_i_0_(cby_9__2__4_right_grid_left_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_f2a_i_0_(cby_9__2__4_right_grid_left_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_f2a_i_0_(cby_9__2__4_right_grid_left_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_f2a_i_0_(cby_9__2__4_right_grid_left_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_8__pin_f2a_i_0_(cby_9__2__4_right_grid_left_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_9__pin_f2a_i_0_(cby_9__2__4_right_grid_left_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_10__pin_f2a_i_0_(cby_9__2__4_right_grid_left_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_11__pin_f2a_i_0_(cby_9__2__4_right_grid_left_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_12__pin_f2a_i_0_(cby_9__2__4_right_grid_left_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_13__pin_f2a_i_0_(cby_9__2__4_right_grid_left_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_14__pin_f2a_i_0_(cby_9__2__4_right_grid_left_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_15__pin_f2a_i_0_(cby_9__2__4_right_grid_left_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_16__pin_f2a_i_0_(cby_9__2__4_right_grid_left_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_17__pin_f2a_i_0_(cby_9__2__4_right_grid_left_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_18__pin_f2a_i_0_(cby_9__2__4_right_grid_left_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_19__pin_f2a_i_0_(cby_9__2__4_right_grid_left_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_0_(cby_9__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_1_(cby_9__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_2_(cby_9__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_3_(cby_9__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_4_(cby_9__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_5_(cby_9__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_6_(cby_9__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_7_(cby_9__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_8_(cby_9__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_9_(cby_9__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_0_(cby_9__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_1_(cby_9__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_2_(cby_9__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_3_(cby_9__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_4_(cby_9__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_5_(cby_9__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_6_(cby_9__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_7_(cby_9__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_8_(cby_9__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_9_(cby_9__2__4_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_0_(cby_9__2__4_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_1_(cby_9__2__4_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_2_(cby_9__2__4_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_3_(cby_9__2__4_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_4_(cby_9__2__4_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_5_(cby_9__2__4_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.ccff_tail(cby_9__2__4_ccff_tail));

	cby_9__2_ cby_9__7_ (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.chany_bottom_in(sb_9__2__4_chany_top_out[0:95]),
		.chany_top_in(sb_9__7__0_chany_bottom_out[0:95]),
		.ccff_head(cbx_2__2__29_ccff_tail),
		.chany_bottom_out(cby_9__2__5_chany_bottom_out[0:95]),
		.chany_top_out(cby_9__2__5_chany_top_out[0:95]),
		.right_grid_left_width_0_height_0_subtile_0__pin_f2a_i_0_(cby_9__2__5_right_grid_left_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_f2a_i_0_(cby_9__2__5_right_grid_left_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_f2a_i_0_(cby_9__2__5_right_grid_left_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_f2a_i_0_(cby_9__2__5_right_grid_left_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_f2a_i_0_(cby_9__2__5_right_grid_left_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_f2a_i_0_(cby_9__2__5_right_grid_left_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_f2a_i_0_(cby_9__2__5_right_grid_left_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_f2a_i_0_(cby_9__2__5_right_grid_left_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_8__pin_f2a_i_0_(cby_9__2__5_right_grid_left_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_9__pin_f2a_i_0_(cby_9__2__5_right_grid_left_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_10__pin_f2a_i_0_(cby_9__2__5_right_grid_left_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_11__pin_f2a_i_0_(cby_9__2__5_right_grid_left_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_12__pin_f2a_i_0_(cby_9__2__5_right_grid_left_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_13__pin_f2a_i_0_(cby_9__2__5_right_grid_left_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_14__pin_f2a_i_0_(cby_9__2__5_right_grid_left_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_15__pin_f2a_i_0_(cby_9__2__5_right_grid_left_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_16__pin_f2a_i_0_(cby_9__2__5_right_grid_left_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_17__pin_f2a_i_0_(cby_9__2__5_right_grid_left_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_18__pin_f2a_i_0_(cby_9__2__5_right_grid_left_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.right_grid_left_width_0_height_0_subtile_19__pin_f2a_i_0_(cby_9__2__5_right_grid_left_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_0_(cby_9__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I2_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_1_(cby_9__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I2_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_2_(cby_9__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I2_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_3_(cby_9__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I2_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_4_(cby_9__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I2_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_5_(cby_9__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I2_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_6_(cby_9__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I2_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_7_(cby_9__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I2_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_8_(cby_9__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I2_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I2_9_(cby_9__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I2_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_0_(cby_9__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I3_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_1_(cby_9__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I3_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_2_(cby_9__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I3_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_3_(cby_9__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I3_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_4_(cby_9__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I3_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_5_(cby_9__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I3_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_6_(cby_9__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I3_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_7_(cby_9__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I3_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_8_(cby_9__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I3_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I3_9_(cby_9__2__5_left_grid_right_width_0_height_0_subtile_0__pin_I3_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_0_(cby_9__2__5_left_grid_right_width_0_height_0_subtile_0__pin_IS_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_1_(cby_9__2__5_left_grid_right_width_0_height_0_subtile_0__pin_IS_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_2_(cby_9__2__5_left_grid_right_width_0_height_0_subtile_0__pin_IS_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_3_(cby_9__2__5_left_grid_right_width_0_height_0_subtile_0__pin_IS_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_4_(cby_9__2__5_left_grid_right_width_0_height_0_subtile_0__pin_IS_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_IS_5_(cby_9__2__5_left_grid_right_width_0_height_0_subtile_0__pin_IS_5_),
		.ccff_tail(cby_9__2__5_ccff_tail));

	direct_interc direct_interc_0_ (
		.in(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_0_out));

	direct_interc direct_interc_1_ (
		.in(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_1_out));

	direct_interc direct_interc_2_ (
		.in(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_2_out));

	direct_interc direct_interc_3_ (
		.in(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_3_out));

	direct_interc direct_interc_4_ (
		.in(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_4_out));

	direct_interc direct_interc_5_ (
		.in(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_5_out));

	direct_interc direct_interc_6_ (
		.in(grid_clb_8_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_6_out));

	direct_interc direct_interc_7_ (
		.in(grid_clb_9_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_7_out));

	direct_interc direct_interc_8_ (
		.in(grid_clb_10_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_8_out));

	direct_interc direct_interc_9_ (
		.in(grid_clb_11_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_9_out));

	direct_interc direct_interc_10_ (
		.in(grid_clb_13_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_10_out));

	direct_interc direct_interc_11_ (
		.in(grid_clb_14_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_11_out));

	direct_interc direct_interc_12_ (
		.in(grid_clb_15_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_12_out));

	direct_interc direct_interc_13_ (
		.in(grid_clb_16_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_13_out));

	direct_interc direct_interc_14_ (
		.in(grid_clb_17_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_14_out));

	direct_interc direct_interc_15_ (
		.in(grid_clb_19_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_15_out));

	direct_interc direct_interc_16_ (
		.in(grid_clb_20_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_16_out));

	direct_interc direct_interc_17_ (
		.in(grid_clb_21_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_17_out));

	direct_interc direct_interc_18_ (
		.in(grid_clb_22_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_18_out));

	direct_interc direct_interc_19_ (
		.in(grid_clb_23_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_19_out));

	direct_interc direct_interc_20_ (
		.in(grid_clb_25_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_20_out));

	direct_interc direct_interc_21_ (
		.in(grid_clb_26_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_21_out));

	direct_interc direct_interc_22_ (
		.in(grid_clb_27_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_22_out));

	direct_interc direct_interc_23_ (
		.in(grid_clb_28_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_23_out));

	direct_interc direct_interc_24_ (
		.in(grid_clb_29_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_24_out));

	direct_interc direct_interc_25_ (
		.in(grid_clb_31_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_25_out));

	direct_interc direct_interc_26_ (
		.in(grid_clb_32_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_26_out));

	direct_interc direct_interc_27_ (
		.in(grid_clb_33_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_27_out));

	direct_interc direct_interc_28_ (
		.in(grid_clb_34_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_28_out));

	direct_interc direct_interc_29_ (
		.in(grid_clb_35_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_29_out));

endmodule
// ----- END Verilog module for fpga_top -----

//----- Default net type -----
`default_nettype none




