//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Fabric Netlist Summary
//	Author: Xifan TANG
//	Organization: University of Utah
//-------------------------------------------
//----- Time scale -----
`timescale 1ns / 1ps

// ------ Include defines: preproc flags -----
`include "../../SRC/fpga_defines.v"
`include "../../SRC/CustomModules/bram/rtl/dti_dp_tm16ffcll_1024x18_t8bw2x_m_hc.v"

`include "/cadlib/gemini/TSMC16NMFFC/library/std_cells/dti/7p5t/rev_220704/220704_dti_tm16ffc_90c_7p5t_stdcells_rev1p0p1_rapid_fe_views_svt/220704_dti_tm16ffc_90c_7p5t_stdcells_rev1p0p1_rapid/verilog/dti_tm16ffc_90c_7p5t_stdcells_rev1p0p0.v"
// ------ Include user-defined netlists -----
`include "../../sim/dti_tm16ffc_90c_7p5t_stdcells_rev1p0p0.v"
`include "../../SRC/CustomModules/QL_PREIO_dti.v"
`include "../../SRC/CustomModules/QL_IOFF_dti.v"
`include "../../SRC/CustomModules/QL_XOR_MUX2_dti.v"
`include "../../SRC/CustomModules/GC_FF_dti.v"
`include "../../SRC/CustomModules/rs_ccff.v"
`include "../../SRC/CustomModules/RS_CCFF_dti.v"
`include "../../SRC/CustomModules/ql_preio.v"
`include "../../SRC/CustomModules/ql_ioff.v"
`include "../../SRC/CustomModules/ql_xor_mux2.v"
`include "../../SRC/CustomModules/ql_ff.v"
`include "../../SRC/CustomModules/gc_ff.v"
`include "../../SRC/CustomModules/ql_dsp.v"
`include "../../SRC/CustomModules/QL_DSP.v"
`include "../../SRC/CustomModules/QL_TDP36K.v"
`include "../../SRC/CustomModules/QL_BRAM.v"
// ------ Include primitive module netlists -----
`include "../../SRC/sub_module/inv_buf_passgate.v"
`include "../../SRC/sub_module/arch_encoder.v"
`include "../../SRC/sub_module/local_encoder.v"
`include "../../SRC/sub_module/mux_primitives.v"
`include "../../SRC/sub_module/muxes.v"
`include "../../SRC/sub_module/luts.v"
`include "../../SRC/sub_module/wires.v"
`include "../../SRC/sub_module/memories.v"
`include "../../SRC/sub_module/shift_register_banks.v"

// ------ Include logic block netlists -----
`include "../../SRC/lb/logical_tile_io_mode_physical__iopad_mode_default__ff.v"
`include "../../SRC/lb/logical_tile_io_mode_physical__iopad_mode_default__pad.v"
`include "../../SRC/lb/logical_tile_io_mode_physical__iopad.v"
`include "../../SRC/lb/logical_tile_io_mode_io_.v"
`include "../../SRC/lb/logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut6.v"
`include "../../SRC/lb/logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__adder_carry.v"
`include "../../SRC/lb/logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic.v"
`include "../../SRC/lb/logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_phy.v"
`include "../../SRC/lb/logical_tile_clb_mode_default__fle_mode_physical__fabric.v"
`include "../../SRC/lb/logical_tile_clb_mode_default__fle.v"
`include "../../SRC/lb/logical_tile_clb_mode_clb_.v"
`include "../../SRC/lb/logical_tile_dsp_mode_physical__dsp_phy.v"
`include "../../SRC/lb/logical_tile_dsp_mode_dsp_.v"
`include "../../SRC/lb/logical_tile_bram_mode_physical__bram_phy.v"
`include "../../SRC/lb/logical_tile_bram_mode_bram_.v"
`include "../../SRC/lb/grid_io_top.v"
`include "../../SRC/lb/grid_io_right.v"
`include "../../SRC/lb/grid_io_bottom.v"
`include "../../SRC/lb/grid_io_left.v"
`include "../../SRC/lb/grid_clb.v"
`include "../../SRC/lb/grid_dsp.v"
`include "../../SRC/lb/grid_bram.v"

// ------ Include routing module netlists -----
`include "../../SRC/routing/sb_0__0_.v"
`include "../../SRC/routing/sb_0__1_.v"
`include "../../SRC/routing/sb_0__8_.v"
`include "../../SRC/routing/sb_1__0_.v"
`include "../../SRC/routing/sb_1__1_.v"
`include "../../SRC/routing/sb_1__2_.v"
`include "../../SRC/routing/sb_1__7_.v"
`include "../../SRC/routing/sb_1__8_.v"
`include "../../SRC/routing/sb_2__0_.v"
`include "../../SRC/routing/sb_2__1_.v"
`include "../../SRC/routing/sb_2__2_.v"
`include "../../SRC/routing/sb_2__7_.v"
`include "../../SRC/routing/sb_2__8_.v"
`include "../../SRC/routing/sb_3__1_.v"
`include "../../SRC/routing/sb_3__2_.v"
`include "../../SRC/routing/sb_3__4_.v"
`include "../../SRC/routing/sb_3__7_.v"
`include "../../SRC/routing/sb_4__1_.v"
`include "../../SRC/routing/sb_4__2_.v"
`include "../../SRC/routing/sb_4__3_.v"
`include "../../SRC/routing/sb_4__4_.v"
`include "../../SRC/routing/sb_4__7_.v"
`include "../../SRC/routing/sb_7__1_.v"
`include "../../SRC/routing/sb_7__2_.v"
`include "../../SRC/routing/sb_7__7_.v"
`include "../../SRC/routing/sb_9__1_.v"
`include "../../SRC/routing/sb_9__2_.v"
`include "../../SRC/routing/sb_9__7_.v"
`include "../../SRC/routing/sb_10__0_.v"
`include "../../SRC/routing/sb_10__1_.v"
`include "../../SRC/routing/sb_10__8_.v"
`include "../../SRC/routing/cbx_1__0_.v"
`include "../../SRC/routing/cbx_2__1_.v"
`include "../../SRC/routing/cbx_2__2_.v"
`include "../../SRC/routing/cbx_2__7_.v"
`include "../../SRC/routing/cbx_4__1_.v"
`include "../../SRC/routing/cbx_4__4_.v"
`include "../../SRC/routing/cbx_4__7_.v"
`include "../../SRC/routing/cbx_7__1_.v"
`include "../../SRC/routing/cby_0__1_.v"
`include "../../SRC/routing/cby_1__1_.v"
`include "../../SRC/routing/cby_2__2_.v"
`include "../../SRC/routing/cby_4__2_.v"
`include "../../SRC/routing/cby_4__3_.v"
`include "../../SRC/routing/cby_4__4_.v"
`include "../../SRC/routing/cby_7__2_.v"
`include "../../SRC/routing/cby_7__3_.v"
`include "../../SRC/routing/cby_7__4_.v"
`include "../../SRC/routing/cby_7__5_.v"
`include "../../SRC/routing/cby_7__6_.v"
`include "../../SRC/routing/cby_7__7_.v"
`include "../../SRC/routing/cby_9__1_.v"
`include "../../SRC/routing/cby_9__2_.v"

// ------ Include fabric top-level netlists -----
`include "../../SRC/fpga_top.v"

