//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for Unique Switch Blocks[0][0]
//	Author: Xifan TANG
//	Organization: University of Utah
//-------------------------------------------
//----- Time scale -----
`timescale 1ns / 1ps

//----- Default net type -----
`default_nettype wire

// ----- Verilog module for sb_0__0_ -----
module sb_0__0_(config_enable,
                prog_clock,
                chany_top_in,
                top_right_grid_left_width_0_height_0_subtile_24__pin_a2f_o_0_,
                top_right_grid_left_width_0_height_0_subtile_25__pin_a2f_o_0_,
                top_right_grid_left_width_0_height_0_subtile_26__pin_a2f_o_0_,
                top_right_grid_left_width_0_height_0_subtile_27__pin_a2f_o_0_,
                top_right_grid_left_width_0_height_0_subtile_28__pin_a2f_o_0_,
                top_right_grid_left_width_0_height_0_subtile_29__pin_a2f_o_0_,
                top_right_grid_left_width_0_height_0_subtile_30__pin_a2f_o_0_,
                top_right_grid_left_width_0_height_0_subtile_31__pin_a2f_o_0_,
                top_right_grid_left_width_0_height_0_subtile_32__pin_a2f_o_0_,
                top_right_grid_left_width_0_height_0_subtile_33__pin_a2f_o_0_,
                top_right_grid_left_width_0_height_0_subtile_34__pin_a2f_o_0_,
                top_right_grid_left_width_0_height_0_subtile_35__pin_a2f_o_0_,
                top_right_grid_left_width_0_height_0_subtile_36__pin_a2f_o_0_,
                top_right_grid_left_width_0_height_0_subtile_37__pin_a2f_o_0_,
                top_right_grid_left_width_0_height_0_subtile_38__pin_a2f_o_0_,
                top_right_grid_left_width_0_height_0_subtile_39__pin_a2f_o_0_,
                top_right_grid_left_width_0_height_0_subtile_40__pin_a2f_o_0_,
                top_right_grid_left_width_0_height_0_subtile_41__pin_a2f_o_0_,
                top_right_grid_left_width_0_height_0_subtile_42__pin_a2f_o_0_,
                top_right_grid_left_width_0_height_0_subtile_43__pin_a2f_o_0_,
                top_right_grid_left_width_0_height_0_subtile_44__pin_a2f_o_0_,
                top_right_grid_left_width_0_height_0_subtile_45__pin_a2f_o_0_,
                top_right_grid_left_width_0_height_0_subtile_46__pin_a2f_o_0_,
                top_right_grid_left_width_0_height_0_subtile_47__pin_a2f_o_0_,
                top_right_grid_left_width_0_height_0_subtile_48__pin_a2f_o_0_,
                top_right_grid_left_width_0_height_0_subtile_49__pin_a2f_o_0_,
                top_right_grid_left_width_0_height_0_subtile_50__pin_a2f_o_0_,
                top_right_grid_left_width_0_height_0_subtile_51__pin_a2f_o_0_,
                top_right_grid_left_width_0_height_0_subtile_52__pin_a2f_o_0_,
                top_right_grid_left_width_0_height_0_subtile_53__pin_a2f_o_0_,
                top_right_grid_left_width_0_height_0_subtile_54__pin_a2f_o_0_,
                top_right_grid_left_width_0_height_0_subtile_55__pin_a2f_o_0_,
                top_right_grid_left_width_0_height_0_subtile_56__pin_a2f_o_0_,
                top_right_grid_left_width_0_height_0_subtile_57__pin_a2f_o_0_,
                top_right_grid_left_width_0_height_0_subtile_58__pin_a2f_o_0_,
                top_right_grid_left_width_0_height_0_subtile_59__pin_a2f_o_0_,
                top_right_grid_left_width_0_height_0_subtile_60__pin_a2f_o_0_,
                top_right_grid_left_width_0_height_0_subtile_61__pin_a2f_o_0_,
                top_right_grid_left_width_0_height_0_subtile_62__pin_a2f_o_0_,
                top_right_grid_left_width_0_height_0_subtile_63__pin_a2f_o_0_,
                top_right_grid_left_width_0_height_0_subtile_64__pin_a2f_o_0_,
                top_right_grid_left_width_0_height_0_subtile_65__pin_a2f_o_0_,
                top_right_grid_left_width_0_height_0_subtile_66__pin_a2f_o_0_,
                top_right_grid_left_width_0_height_0_subtile_67__pin_a2f_o_0_,
                top_right_grid_left_width_0_height_0_subtile_68__pin_a2f_o_0_,
                top_right_grid_left_width_0_height_0_subtile_69__pin_a2f_o_0_,
                top_right_grid_left_width_0_height_0_subtile_70__pin_a2f_o_0_,
                top_right_grid_left_width_0_height_0_subtile_71__pin_a2f_o_0_,
                chanx_right_in,
                ccff_head,
                chany_top_out,
                chanx_right_out,
                ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_clock;
//----- INPUT PORTS -----
input [0:95] chany_top_in;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_24__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_25__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_26__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_27__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_28__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_29__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_30__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_31__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_32__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_33__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_34__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_35__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_36__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_37__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_38__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_39__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_40__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_41__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_42__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_43__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_44__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_45__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_46__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_47__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_48__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_49__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_50__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_51__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_52__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_53__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_54__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_55__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_56__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_57__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_58__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_59__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_60__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_61__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_62__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_63__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_64__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_65__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_66__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_67__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_68__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_69__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_70__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_71__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:95] chanx_right_in;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:95] chany_top_out;
//----- OUTPUT PORTS -----
output [0:95] chanx_right_out;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:1] mux_tree_tapbuf_L2SB_size3_0_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size3_0_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size3_1_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size3_1_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size3_2_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size3_2_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size3_3_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size3_3_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size3_4_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size3_4_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size3_5_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size3_5_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size3_6_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size3_6_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size3_7_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size3_7_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size3_8_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size3_8_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_0_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_0_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_1_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_1_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_2_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_2_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_3_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_3_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_4_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_4_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_5_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_5_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_6_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_6_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_7_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_7_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_8_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_8_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_9_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_9_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_0_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_0_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_10_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_10_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_1_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_1_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_2_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_2_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_3_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_3_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_4_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_4_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_5_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_5_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_6_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_6_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_7_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_7_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_8_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_8_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_9_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_9_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_0_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_0_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_10_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_10_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_11_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_11_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_12_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_12_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_13_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_13_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_14_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_14_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_15_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_15_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_16_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_16_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_17_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_17_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_18_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_18_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_19_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_19_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_1_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_1_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_20_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_20_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_21_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_21_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_22_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_22_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_23_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_23_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_24_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_24_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_25_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_25_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_26_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_26_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_27_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_27_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_28_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_28_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_29_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_29_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_2_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_2_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_30_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_30_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_31_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_31_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_32_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_32_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_33_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_33_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_34_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_34_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_35_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_35_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_36_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_36_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_37_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_37_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_38_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_38_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_39_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_39_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_3_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_3_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_40_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_40_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_41_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_41_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_42_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_42_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_43_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_43_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_44_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_44_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_45_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_45_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_46_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_46_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_47_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_47_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_48_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_48_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_49_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_49_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_4_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_4_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_50_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_50_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_51_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_51_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_52_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_52_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_53_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_53_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_54_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_54_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_55_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_55_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_56_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_56_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_57_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_57_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_58_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_58_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_59_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_59_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_5_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_5_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_60_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_60_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_61_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_61_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_62_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_62_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_63_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_63_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_64_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_64_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_65_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_65_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_6_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_6_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_7_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_7_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_8_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_8_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_9_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_9_sram_inv;

// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[1] = chany_top_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[2] = chany_top_in[1];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[3] = chany_top_in[2];
// ----- Local connection due to Wire 3 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[4] = chany_top_in[3];
// ----- Local connection due to Wire 4 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[5] = chany_top_in[4];
// ----- Local connection due to Wire 5 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[6] = chany_top_in[5];
// ----- Local connection due to Wire 6 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[7] = chany_top_in[6];
// ----- Local connection due to Wire 7 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[8] = chany_top_in[7];
// ----- Local connection due to Wire 8 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[9] = chany_top_in[8];
// ----- Local connection due to Wire 9 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[10] = chany_top_in[9];
// ----- Local connection due to Wire 10 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[11] = chany_top_in[10];
// ----- Local connection due to Wire 11 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[12] = chany_top_in[11];
// ----- Local connection due to Wire 12 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[13] = chany_top_in[12];
// ----- Local connection due to Wire 13 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[14] = chany_top_in[13];
// ----- Local connection due to Wire 14 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[15] = chany_top_in[14];
// ----- Local connection due to Wire 15 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[16] = chany_top_in[15];
// ----- Local connection due to Wire 16 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[17] = chany_top_in[16];
// ----- Local connection due to Wire 17 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[18] = chany_top_in[17];
// ----- Local connection due to Wire 18 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[19] = chany_top_in[18];
// ----- Local connection due to Wire 19 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[20] = chany_top_in[19];
// ----- Local connection due to Wire 20 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[21] = chany_top_in[20];
// ----- Local connection due to Wire 21 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[22] = chany_top_in[21];
// ----- Local connection due to Wire 22 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[23] = chany_top_in[22];
// ----- Local connection due to Wire 23 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[24] = chany_top_in[23];
// ----- Local connection due to Wire 24 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[25] = chany_top_in[24];
// ----- Local connection due to Wire 25 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[26] = chany_top_in[25];
// ----- Local connection due to Wire 26 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[27] = chany_top_in[26];
// ----- Local connection due to Wire 27 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[28] = chany_top_in[27];
// ----- Local connection due to Wire 28 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[29] = chany_top_in[28];
// ----- Local connection due to Wire 29 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[30] = chany_top_in[29];
// ----- Local connection due to Wire 30 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[31] = chany_top_in[30];
// ----- Local connection due to Wire 31 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[32] = chany_top_in[31];
// ----- Local connection due to Wire 32 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[33] = chany_top_in[32];
// ----- Local connection due to Wire 33 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[34] = chany_top_in[33];
// ----- Local connection due to Wire 34 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[35] = chany_top_in[34];
// ----- Local connection due to Wire 35 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[36] = chany_top_in[35];
// ----- Local connection due to Wire 36 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[37] = chany_top_in[36];
// ----- Local connection due to Wire 37 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[38] = chany_top_in[37];
// ----- Local connection due to Wire 38 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[39] = chany_top_in[38];
// ----- Local connection due to Wire 39 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[40] = chany_top_in[39];
// ----- Local connection due to Wire 40 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[41] = chany_top_in[40];
// ----- Local connection due to Wire 41 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[42] = chany_top_in[41];
// ----- Local connection due to Wire 42 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[43] = chany_top_in[42];
// ----- Local connection due to Wire 43 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[44] = chany_top_in[43];
// ----- Local connection due to Wire 44 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[45] = chany_top_in[44];
// ----- Local connection due to Wire 45 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[46] = chany_top_in[45];
// ----- Local connection due to Wire 46 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[47] = chany_top_in[46];
// ----- Local connection due to Wire 47 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[48] = chany_top_in[47];
// ----- Local connection due to Wire 48 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[49] = chany_top_in[48];
// ----- Local connection due to Wire 49 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[50] = chany_top_in[49];
// ----- Local connection due to Wire 50 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[51] = chany_top_in[50];
// ----- Local connection due to Wire 51 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[52] = chany_top_in[51];
// ----- Local connection due to Wire 52 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[53] = chany_top_in[52];
// ----- Local connection due to Wire 53 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[54] = chany_top_in[53];
// ----- Local connection due to Wire 54 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[55] = chany_top_in[54];
// ----- Local connection due to Wire 55 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[56] = chany_top_in[55];
// ----- Local connection due to Wire 56 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[57] = chany_top_in[56];
// ----- Local connection due to Wire 57 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[58] = chany_top_in[57];
// ----- Local connection due to Wire 58 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[59] = chany_top_in[58];
// ----- Local connection due to Wire 59 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[60] = chany_top_in[59];
// ----- Local connection due to Wire 60 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[61] = chany_top_in[60];
// ----- Local connection due to Wire 61 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[62] = chany_top_in[61];
// ----- Local connection due to Wire 62 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[63] = chany_top_in[62];
// ----- Local connection due to Wire 63 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[64] = chany_top_in[63];
// ----- Local connection due to Wire 64 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[65] = chany_top_in[64];
// ----- Local connection due to Wire 65 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[66] = chany_top_in[65];
// ----- Local connection due to Wire 66 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[67] = chany_top_in[66];
// ----- Local connection due to Wire 67 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[68] = chany_top_in[67];
// ----- Local connection due to Wire 68 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[69] = chany_top_in[68];
// ----- Local connection due to Wire 69 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[70] = chany_top_in[69];
// ----- Local connection due to Wire 70 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[71] = chany_top_in[70];
// ----- Local connection due to Wire 71 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[72] = chany_top_in[71];
// ----- Local connection due to Wire 72 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[73] = chany_top_in[72];
// ----- Local connection due to Wire 73 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[74] = chany_top_in[73];
// ----- Local connection due to Wire 74 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[75] = chany_top_in[74];
// ----- Local connection due to Wire 75 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[76] = chany_top_in[75];
// ----- Local connection due to Wire 76 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[77] = chany_top_in[76];
// ----- Local connection due to Wire 77 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[78] = chany_top_in[77];
// ----- Local connection due to Wire 78 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[79] = chany_top_in[78];
// ----- Local connection due to Wire 79 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[80] = chany_top_in[79];
// ----- Local connection due to Wire 80 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[81] = chany_top_in[80];
// ----- Local connection due to Wire 81 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[82] = chany_top_in[81];
// ----- Local connection due to Wire 82 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[83] = chany_top_in[82];
// ----- Local connection due to Wire 83 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[84] = chany_top_in[83];
// ----- Local connection due to Wire 84 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[85] = chany_top_in[84];
// ----- Local connection due to Wire 85 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[86] = chany_top_in[85];
// ----- Local connection due to Wire 86 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[87] = chany_top_in[86];
// ----- Local connection due to Wire 87 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[88] = chany_top_in[87];
// ----- Local connection due to Wire 88 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[89] = chany_top_in[88];
// ----- Local connection due to Wire 89 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[90] = chany_top_in[89];
// ----- Local connection due to Wire 90 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[91] = chany_top_in[90];
// ----- Local connection due to Wire 91 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[92] = chany_top_in[91];
// ----- Local connection due to Wire 92 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[93] = chany_top_in[92];
// ----- Local connection due to Wire 93 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[94] = chany_top_in[93];
// ----- Local connection due to Wire 94 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[95] = chany_top_in[94];
// ----- Local connection due to Wire 95 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[0] = chany_top_in[95];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	mux_tree_tapbuf_L2SB_size4 mux_top_track_0 (
		.in({top_right_grid_left_width_0_height_0_subtile_24__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_43__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_62__pin_a2f_o_0_, chanx_right_in[1]}),
		.sram(mux_tree_tapbuf_L2SB_size4_0_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_0_sram_inv[0:1]),
		.out(chany_top_out[0]));

	mux_tree_tapbuf_L2SB_size4 mux_top_track_2 (
		.in({top_right_grid_left_width_0_height_0_subtile_25__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_44__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_63__pin_a2f_o_0_, chanx_right_in[2]}),
		.sram(mux_tree_tapbuf_L2SB_size4_1_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_1_sram_inv[0:1]),
		.out(chany_top_out[1]));

	mux_tree_tapbuf_L2SB_size4 mux_top_track_4 (
		.in({top_right_grid_left_width_0_height_0_subtile_26__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_45__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_64__pin_a2f_o_0_, chanx_right_in[3]}),
		.sram(mux_tree_tapbuf_L2SB_size4_2_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_2_sram_inv[0:1]),
		.out(chany_top_out[2]));

	mux_tree_tapbuf_L2SB_size4 mux_top_track_6 (
		.in({top_right_grid_left_width_0_height_0_subtile_27__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_46__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_65__pin_a2f_o_0_, chanx_right_in[4]}),
		.sram(mux_tree_tapbuf_L2SB_size4_3_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_3_sram_inv[0:1]),
		.out(chany_top_out[3]));

	mux_tree_tapbuf_L2SB_size4 mux_top_track_8 (
		.in({top_right_grid_left_width_0_height_0_subtile_28__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_47__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_66__pin_a2f_o_0_, chanx_right_in[5]}),
		.sram(mux_tree_tapbuf_L2SB_size4_4_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_4_sram_inv[0:1]),
		.out(chany_top_out[4]));

	mux_tree_tapbuf_L2SB_size4 mux_top_track_10 (
		.in({top_right_grid_left_width_0_height_0_subtile_29__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_48__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_67__pin_a2f_o_0_, chanx_right_in[6]}),
		.sram(mux_tree_tapbuf_L2SB_size4_5_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_5_sram_inv[0:1]),
		.out(chany_top_out[5]));

	mux_tree_tapbuf_L2SB_size4 mux_top_track_12 (
		.in({top_right_grid_left_width_0_height_0_subtile_30__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_49__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_68__pin_a2f_o_0_, chanx_right_in[7]}),
		.sram(mux_tree_tapbuf_L2SB_size4_6_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_6_sram_inv[0:1]),
		.out(chany_top_out[6]));

	mux_tree_tapbuf_L2SB_size4 mux_top_track_14 (
		.in({top_right_grid_left_width_0_height_0_subtile_31__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_50__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_69__pin_a2f_o_0_, chanx_right_in[8]}),
		.sram(mux_tree_tapbuf_L2SB_size4_7_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_7_sram_inv[0:1]),
		.out(chany_top_out[7]));

	mux_tree_tapbuf_L2SB_size4 mux_top_track_16 (
		.in({top_right_grid_left_width_0_height_0_subtile_32__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_51__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_70__pin_a2f_o_0_, chanx_right_in[9]}),
		.sram(mux_tree_tapbuf_L2SB_size4_8_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_8_sram_inv[0:1]),
		.out(chany_top_out[8]));

	mux_tree_tapbuf_L2SB_size4 mux_top_track_18 (
		.in({top_right_grid_left_width_0_height_0_subtile_33__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_52__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_71__pin_a2f_o_0_, chanx_right_in[10]}),
		.sram(mux_tree_tapbuf_L2SB_size4_9_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_9_sram_inv[0:1]),
		.out(chany_top_out[9]));

	mux_tree_tapbuf_L2SB_size4_mem mem_top_track_0 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(ccff_head),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_0_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_0_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_top_track_2 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_1_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_1_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_top_track_4 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_2_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_2_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_top_track_6 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_3_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_3_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_top_track_8 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_4_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_4_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_top_track_10 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_5_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_5_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_top_track_12 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_6_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_6_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_top_track_14 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_7_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_7_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_top_track_16 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_8_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_8_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_top_track_18 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_9_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_9_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size3 mux_top_track_20 (
		.in({top_right_grid_left_width_0_height_0_subtile_34__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_53__pin_a2f_o_0_, chanx_right_in[11]}),
		.sram(mux_tree_tapbuf_L2SB_size3_0_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size3_0_sram_inv[0:1]),
		.out(chany_top_out[10]));

	mux_tree_tapbuf_L2SB_size3 mux_top_track_22 (
		.in({top_right_grid_left_width_0_height_0_subtile_35__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_54__pin_a2f_o_0_, chanx_right_in[12]}),
		.sram(mux_tree_tapbuf_L2SB_size3_1_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size3_1_sram_inv[0:1]),
		.out(chany_top_out[11]));

	mux_tree_tapbuf_L2SB_size3 mux_top_track_24 (
		.in({top_right_grid_left_width_0_height_0_subtile_36__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_55__pin_a2f_o_0_, chanx_right_in[13]}),
		.sram(mux_tree_tapbuf_L2SB_size3_2_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size3_2_sram_inv[0:1]),
		.out(chany_top_out[12]));

	mux_tree_tapbuf_L2SB_size3 mux_top_track_26 (
		.in({top_right_grid_left_width_0_height_0_subtile_37__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_56__pin_a2f_o_0_, chanx_right_in[14]}),
		.sram(mux_tree_tapbuf_L2SB_size3_3_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size3_3_sram_inv[0:1]),
		.out(chany_top_out[13]));

	mux_tree_tapbuf_L2SB_size3 mux_top_track_28 (
		.in({top_right_grid_left_width_0_height_0_subtile_38__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_57__pin_a2f_o_0_, chanx_right_in[15]}),
		.sram(mux_tree_tapbuf_L2SB_size3_4_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size3_4_sram_inv[0:1]),
		.out(chany_top_out[14]));

	mux_tree_tapbuf_L2SB_size3 mux_top_track_30 (
		.in({top_right_grid_left_width_0_height_0_subtile_39__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_58__pin_a2f_o_0_, chanx_right_in[16]}),
		.sram(mux_tree_tapbuf_L2SB_size3_5_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size3_5_sram_inv[0:1]),
		.out(chany_top_out[15]));

	mux_tree_tapbuf_L2SB_size3 mux_top_track_32 (
		.in({top_right_grid_left_width_0_height_0_subtile_40__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_59__pin_a2f_o_0_, chanx_right_in[17]}),
		.sram(mux_tree_tapbuf_L2SB_size3_6_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size3_6_sram_inv[0:1]),
		.out(chany_top_out[16]));

	mux_tree_tapbuf_L2SB_size3 mux_top_track_34 (
		.in({top_right_grid_left_width_0_height_0_subtile_41__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_60__pin_a2f_o_0_, chanx_right_in[18]}),
		.sram(mux_tree_tapbuf_L2SB_size3_7_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size3_7_sram_inv[0:1]),
		.out(chany_top_out[17]));

	mux_tree_tapbuf_L2SB_size3 mux_top_track_36 (
		.in({top_right_grid_left_width_0_height_0_subtile_42__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_61__pin_a2f_o_0_, chanx_right_in[19]}),
		.sram(mux_tree_tapbuf_L2SB_size3_8_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size3_8_sram_inv[0:1]),
		.out(chany_top_out[18]));

	mux_tree_tapbuf_L2SB_size3_mem mem_top_track_20 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size3_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size3_0_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size3_0_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size3_mem mem_top_track_22 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size3_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size3_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size3_1_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size3_1_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size3_mem mem_top_track_24 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size3_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size3_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size3_2_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size3_2_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size3_mem mem_top_track_26 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size3_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size3_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size3_3_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size3_3_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size3_mem mem_top_track_28 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size3_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size3_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size3_4_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size3_4_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size3_mem mem_top_track_30 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size3_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size3_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size3_5_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size3_5_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size3_mem mem_top_track_32 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size3_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size3_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size3_6_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size3_6_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size3_mem mem_top_track_34 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size3_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size3_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size3_7_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size3_7_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size3_mem mem_top_track_36 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size3_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size3_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size3_8_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size3_8_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_38 (
		.in({top_right_grid_left_width_0_height_0_subtile_24__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_31__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_38__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_45__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_52__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_59__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_66__pin_a2f_o_0_, chanx_right_in[20]}),
		.sram(mux_tree_tapbuf_L4SB_size8_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_0_sram_inv[0:2]),
		.out(chany_top_out[19]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_40 (
		.in({top_right_grid_left_width_0_height_0_subtile_25__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_32__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_39__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_46__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_53__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_60__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_67__pin_a2f_o_0_, chanx_right_in[21]}),
		.sram(mux_tree_tapbuf_L4SB_size8_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_1_sram_inv[0:2]),
		.out(chany_top_out[20]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_42 (
		.in({top_right_grid_left_width_0_height_0_subtile_26__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_33__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_40__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_47__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_54__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_61__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_68__pin_a2f_o_0_, chanx_right_in[22]}),
		.sram(mux_tree_tapbuf_L4SB_size8_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_2_sram_inv[0:2]),
		.out(chany_top_out[21]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_44 (
		.in({top_right_grid_left_width_0_height_0_subtile_27__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_34__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_41__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_48__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_55__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_62__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_69__pin_a2f_o_0_, chanx_right_in[23]}),
		.sram(mux_tree_tapbuf_L4SB_size8_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_3_sram_inv[0:2]),
		.out(chany_top_out[22]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_46 (
		.in({top_right_grid_left_width_0_height_0_subtile_28__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_35__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_42__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_49__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_56__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_63__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_70__pin_a2f_o_0_, chanx_right_in[24]}),
		.sram(mux_tree_tapbuf_L4SB_size8_4_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_4_sram_inv[0:2]),
		.out(chany_top_out[23]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_48 (
		.in({top_right_grid_left_width_0_height_0_subtile_29__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_36__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_43__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_50__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_57__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_64__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_71__pin_a2f_o_0_, chanx_right_in[25]}),
		.sram(mux_tree_tapbuf_L4SB_size8_5_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_5_sram_inv[0:2]),
		.out(chany_top_out[24]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_52 (
		.in({top_right_grid_left_width_0_height_0_subtile_24__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_31__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_38__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_45__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_52__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_59__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_66__pin_a2f_o_0_, chanx_right_in[27]}),
		.sram(mux_tree_tapbuf_L4SB_size8_6_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_6_sram_inv[0:2]),
		.out(chany_top_out[26]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_54 (
		.in({top_right_grid_left_width_0_height_0_subtile_25__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_32__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_39__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_46__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_53__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_60__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_67__pin_a2f_o_0_, chanx_right_in[28]}),
		.sram(mux_tree_tapbuf_L4SB_size8_7_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_7_sram_inv[0:2]),
		.out(chany_top_out[27]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_56 (
		.in({top_right_grid_left_width_0_height_0_subtile_26__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_33__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_40__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_47__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_54__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_61__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_68__pin_a2f_o_0_, chanx_right_in[29]}),
		.sram(mux_tree_tapbuf_L4SB_size8_8_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_8_sram_inv[0:2]),
		.out(chany_top_out[28]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_58 (
		.in({top_right_grid_left_width_0_height_0_subtile_27__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_34__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_41__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_48__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_55__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_62__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_69__pin_a2f_o_0_, chanx_right_in[30]}),
		.sram(mux_tree_tapbuf_L4SB_size8_9_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_9_sram_inv[0:2]),
		.out(chany_top_out[29]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_60 (
		.in({top_right_grid_left_width_0_height_0_subtile_28__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_35__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_42__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_49__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_56__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_63__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_70__pin_a2f_o_0_, chanx_right_in[31]}),
		.sram(mux_tree_tapbuf_L4SB_size8_10_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_10_sram_inv[0:2]),
		.out(chany_top_out[30]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_62 (
		.in({top_right_grid_left_width_0_height_0_subtile_29__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_36__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_43__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_50__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_57__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_64__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_71__pin_a2f_o_0_, chanx_right_in[32]}),
		.sram(mux_tree_tapbuf_L4SB_size8_11_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_11_sram_inv[0:2]),
		.out(chany_top_out[31]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_66 (
		.in({top_right_grid_left_width_0_height_0_subtile_24__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_31__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_38__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_45__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_52__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_59__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_66__pin_a2f_o_0_, chanx_right_in[34]}),
		.sram(mux_tree_tapbuf_L4SB_size8_12_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_12_sram_inv[0:2]),
		.out(chany_top_out[33]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_68 (
		.in({top_right_grid_left_width_0_height_0_subtile_25__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_32__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_39__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_46__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_53__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_60__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_67__pin_a2f_o_0_, chanx_right_in[35]}),
		.sram(mux_tree_tapbuf_L4SB_size8_13_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_13_sram_inv[0:2]),
		.out(chany_top_out[34]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_70 (
		.in({top_right_grid_left_width_0_height_0_subtile_26__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_33__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_40__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_47__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_54__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_61__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_68__pin_a2f_o_0_, chanx_right_in[36]}),
		.sram(mux_tree_tapbuf_L4SB_size8_14_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_14_sram_inv[0:2]),
		.out(chany_top_out[35]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_72 (
		.in({top_right_grid_left_width_0_height_0_subtile_27__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_34__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_41__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_48__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_55__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_62__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_69__pin_a2f_o_0_, chanx_right_in[37]}),
		.sram(mux_tree_tapbuf_L4SB_size8_15_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_15_sram_inv[0:2]),
		.out(chany_top_out[36]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_74 (
		.in({top_right_grid_left_width_0_height_0_subtile_28__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_35__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_42__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_49__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_56__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_63__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_70__pin_a2f_o_0_, chanx_right_in[38]}),
		.sram(mux_tree_tapbuf_L4SB_size8_16_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_16_sram_inv[0:2]),
		.out(chany_top_out[37]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_76 (
		.in({top_right_grid_left_width_0_height_0_subtile_29__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_36__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_43__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_50__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_57__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_64__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_71__pin_a2f_o_0_, chanx_right_in[39]}),
		.sram(mux_tree_tapbuf_L4SB_size8_17_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_17_sram_inv[0:2]),
		.out(chany_top_out[38]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_80 (
		.in({top_right_grid_left_width_0_height_0_subtile_24__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_31__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_38__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_45__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_52__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_59__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_66__pin_a2f_o_0_, chanx_right_in[41]}),
		.sram(mux_tree_tapbuf_L4SB_size8_18_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_18_sram_inv[0:2]),
		.out(chany_top_out[40]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_82 (
		.in({top_right_grid_left_width_0_height_0_subtile_25__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_32__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_39__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_46__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_53__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_60__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_67__pin_a2f_o_0_, chanx_right_in[42]}),
		.sram(mux_tree_tapbuf_L4SB_size8_19_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_19_sram_inv[0:2]),
		.out(chany_top_out[41]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_84 (
		.in({top_right_grid_left_width_0_height_0_subtile_26__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_33__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_40__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_47__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_54__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_61__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_68__pin_a2f_o_0_, chanx_right_in[43]}),
		.sram(mux_tree_tapbuf_L4SB_size8_20_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_20_sram_inv[0:2]),
		.out(chany_top_out[42]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_86 (
		.in({top_right_grid_left_width_0_height_0_subtile_27__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_34__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_41__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_48__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_55__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_62__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_69__pin_a2f_o_0_, chanx_right_in[44]}),
		.sram(mux_tree_tapbuf_L4SB_size8_21_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_21_sram_inv[0:2]),
		.out(chany_top_out[43]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_88 (
		.in({top_right_grid_left_width_0_height_0_subtile_28__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_35__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_42__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_49__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_56__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_63__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_70__pin_a2f_o_0_, chanx_right_in[45]}),
		.sram(mux_tree_tapbuf_L4SB_size8_22_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_22_sram_inv[0:2]),
		.out(chany_top_out[44]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_90 (
		.in({top_right_grid_left_width_0_height_0_subtile_29__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_36__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_43__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_50__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_57__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_64__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_71__pin_a2f_o_0_, chanx_right_in[46]}),
		.sram(mux_tree_tapbuf_L4SB_size8_23_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_23_sram_inv[0:2]),
		.out(chany_top_out[45]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_94 (
		.in({top_right_grid_left_width_0_height_0_subtile_24__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_31__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_38__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_45__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_52__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_59__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_66__pin_a2f_o_0_, chanx_right_in[48]}),
		.sram(mux_tree_tapbuf_L4SB_size8_24_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_24_sram_inv[0:2]),
		.out(chany_top_out[47]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_96 (
		.in({top_right_grid_left_width_0_height_0_subtile_25__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_32__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_39__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_46__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_53__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_60__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_67__pin_a2f_o_0_, chanx_right_in[49]}),
		.sram(mux_tree_tapbuf_L4SB_size8_25_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_25_sram_inv[0:2]),
		.out(chany_top_out[48]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_98 (
		.in({top_right_grid_left_width_0_height_0_subtile_26__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_33__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_40__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_47__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_54__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_61__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_68__pin_a2f_o_0_, chanx_right_in[50]}),
		.sram(mux_tree_tapbuf_L4SB_size8_26_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_26_sram_inv[0:2]),
		.out(chany_top_out[49]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_100 (
		.in({top_right_grid_left_width_0_height_0_subtile_27__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_34__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_41__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_48__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_55__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_62__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_69__pin_a2f_o_0_, chanx_right_in[51]}),
		.sram(mux_tree_tapbuf_L4SB_size8_27_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_27_sram_inv[0:2]),
		.out(chany_top_out[50]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_102 (
		.in({top_right_grid_left_width_0_height_0_subtile_28__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_35__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_42__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_49__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_56__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_63__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_70__pin_a2f_o_0_, chanx_right_in[52]}),
		.sram(mux_tree_tapbuf_L4SB_size8_28_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_28_sram_inv[0:2]),
		.out(chany_top_out[51]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_104 (
		.in({top_right_grid_left_width_0_height_0_subtile_29__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_36__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_43__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_50__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_57__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_64__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_71__pin_a2f_o_0_, chanx_right_in[53]}),
		.sram(mux_tree_tapbuf_L4SB_size8_29_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_29_sram_inv[0:2]),
		.out(chany_top_out[52]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_108 (
		.in({top_right_grid_left_width_0_height_0_subtile_24__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_31__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_38__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_45__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_52__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_59__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_66__pin_a2f_o_0_, chanx_right_in[55]}),
		.sram(mux_tree_tapbuf_L4SB_size8_30_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_30_sram_inv[0:2]),
		.out(chany_top_out[54]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_110 (
		.in({top_right_grid_left_width_0_height_0_subtile_25__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_32__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_39__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_46__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_53__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_60__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_67__pin_a2f_o_0_, chanx_right_in[56]}),
		.sram(mux_tree_tapbuf_L4SB_size8_31_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_31_sram_inv[0:2]),
		.out(chany_top_out[55]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_112 (
		.in({top_right_grid_left_width_0_height_0_subtile_26__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_33__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_40__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_47__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_54__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_61__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_68__pin_a2f_o_0_, chanx_right_in[57]}),
		.sram(mux_tree_tapbuf_L4SB_size8_32_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_32_sram_inv[0:2]),
		.out(chany_top_out[56]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_114 (
		.in({top_right_grid_left_width_0_height_0_subtile_27__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_34__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_41__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_48__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_55__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_62__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_69__pin_a2f_o_0_, chanx_right_in[58]}),
		.sram(mux_tree_tapbuf_L4SB_size8_33_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_33_sram_inv[0:2]),
		.out(chany_top_out[57]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_116 (
		.in({top_right_grid_left_width_0_height_0_subtile_28__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_35__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_42__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_49__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_56__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_63__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_70__pin_a2f_o_0_, chanx_right_in[59]}),
		.sram(mux_tree_tapbuf_L4SB_size8_34_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_34_sram_inv[0:2]),
		.out(chany_top_out[58]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_118 (
		.in({top_right_grid_left_width_0_height_0_subtile_29__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_36__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_43__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_50__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_57__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_64__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_71__pin_a2f_o_0_, chanx_right_in[60]}),
		.sram(mux_tree_tapbuf_L4SB_size8_35_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_35_sram_inv[0:2]),
		.out(chany_top_out[59]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_122 (
		.in({top_right_grid_left_width_0_height_0_subtile_24__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_31__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_38__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_45__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_52__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_59__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_66__pin_a2f_o_0_, chanx_right_in[62]}),
		.sram(mux_tree_tapbuf_L4SB_size8_36_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_36_sram_inv[0:2]),
		.out(chany_top_out[61]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_124 (
		.in({top_right_grid_left_width_0_height_0_subtile_25__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_32__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_39__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_46__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_53__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_60__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_67__pin_a2f_o_0_, chanx_right_in[63]}),
		.sram(mux_tree_tapbuf_L4SB_size8_37_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_37_sram_inv[0:2]),
		.out(chany_top_out[62]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_126 (
		.in({top_right_grid_left_width_0_height_0_subtile_26__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_33__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_40__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_47__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_54__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_61__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_68__pin_a2f_o_0_, chanx_right_in[64]}),
		.sram(mux_tree_tapbuf_L4SB_size8_38_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_38_sram_inv[0:2]),
		.out(chany_top_out[63]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_128 (
		.in({top_right_grid_left_width_0_height_0_subtile_27__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_34__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_41__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_48__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_55__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_62__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_69__pin_a2f_o_0_, chanx_right_in[65]}),
		.sram(mux_tree_tapbuf_L4SB_size8_39_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_39_sram_inv[0:2]),
		.out(chany_top_out[64]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_130 (
		.in({top_right_grid_left_width_0_height_0_subtile_28__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_35__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_42__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_49__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_56__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_63__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_70__pin_a2f_o_0_, chanx_right_in[66]}),
		.sram(mux_tree_tapbuf_L4SB_size8_40_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_40_sram_inv[0:2]),
		.out(chany_top_out[65]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_132 (
		.in({top_right_grid_left_width_0_height_0_subtile_29__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_36__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_43__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_50__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_57__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_64__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_71__pin_a2f_o_0_, chanx_right_in[67]}),
		.sram(mux_tree_tapbuf_L4SB_size8_41_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_41_sram_inv[0:2]),
		.out(chany_top_out[66]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_136 (
		.in({top_right_grid_left_width_0_height_0_subtile_24__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_31__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_38__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_45__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_52__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_59__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_66__pin_a2f_o_0_, chanx_right_in[69]}),
		.sram(mux_tree_tapbuf_L4SB_size8_42_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_42_sram_inv[0:2]),
		.out(chany_top_out[68]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_138 (
		.in({top_right_grid_left_width_0_height_0_subtile_25__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_32__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_39__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_46__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_53__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_60__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_67__pin_a2f_o_0_, chanx_right_in[70]}),
		.sram(mux_tree_tapbuf_L4SB_size8_43_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_43_sram_inv[0:2]),
		.out(chany_top_out[69]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_140 (
		.in({top_right_grid_left_width_0_height_0_subtile_26__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_33__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_40__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_47__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_54__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_61__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_68__pin_a2f_o_0_, chanx_right_in[71]}),
		.sram(mux_tree_tapbuf_L4SB_size8_44_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_44_sram_inv[0:2]),
		.out(chany_top_out[70]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_142 (
		.in({top_right_grid_left_width_0_height_0_subtile_27__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_34__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_41__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_48__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_55__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_62__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_69__pin_a2f_o_0_, chanx_right_in[72]}),
		.sram(mux_tree_tapbuf_L4SB_size8_45_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_45_sram_inv[0:2]),
		.out(chany_top_out[71]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_144 (
		.in({top_right_grid_left_width_0_height_0_subtile_28__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_35__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_42__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_49__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_56__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_63__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_70__pin_a2f_o_0_, chanx_right_in[73]}),
		.sram(mux_tree_tapbuf_L4SB_size8_46_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_46_sram_inv[0:2]),
		.out(chany_top_out[72]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_146 (
		.in({top_right_grid_left_width_0_height_0_subtile_29__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_36__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_43__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_50__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_57__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_64__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_71__pin_a2f_o_0_, chanx_right_in[74]}),
		.sram(mux_tree_tapbuf_L4SB_size8_47_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_47_sram_inv[0:2]),
		.out(chany_top_out[73]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_150 (
		.in({top_right_grid_left_width_0_height_0_subtile_24__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_31__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_38__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_45__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_52__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_59__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_66__pin_a2f_o_0_, chanx_right_in[76]}),
		.sram(mux_tree_tapbuf_L4SB_size8_48_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_48_sram_inv[0:2]),
		.out(chany_top_out[75]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_152 (
		.in({top_right_grid_left_width_0_height_0_subtile_25__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_32__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_39__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_46__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_53__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_60__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_67__pin_a2f_o_0_, chanx_right_in[77]}),
		.sram(mux_tree_tapbuf_L4SB_size8_49_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_49_sram_inv[0:2]),
		.out(chany_top_out[76]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_154 (
		.in({top_right_grid_left_width_0_height_0_subtile_26__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_33__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_40__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_47__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_54__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_61__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_68__pin_a2f_o_0_, chanx_right_in[78]}),
		.sram(mux_tree_tapbuf_L4SB_size8_50_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_50_sram_inv[0:2]),
		.out(chany_top_out[77]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_156 (
		.in({top_right_grid_left_width_0_height_0_subtile_27__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_34__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_41__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_48__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_55__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_62__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_69__pin_a2f_o_0_, chanx_right_in[79]}),
		.sram(mux_tree_tapbuf_L4SB_size8_51_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_51_sram_inv[0:2]),
		.out(chany_top_out[78]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_158 (
		.in({top_right_grid_left_width_0_height_0_subtile_28__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_35__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_42__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_49__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_56__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_63__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_70__pin_a2f_o_0_, chanx_right_in[80]}),
		.sram(mux_tree_tapbuf_L4SB_size8_52_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_52_sram_inv[0:2]),
		.out(chany_top_out[79]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_160 (
		.in({top_right_grid_left_width_0_height_0_subtile_29__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_36__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_43__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_50__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_57__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_64__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_71__pin_a2f_o_0_, chanx_right_in[81]}),
		.sram(mux_tree_tapbuf_L4SB_size8_53_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_53_sram_inv[0:2]),
		.out(chany_top_out[80]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_164 (
		.in({top_right_grid_left_width_0_height_0_subtile_24__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_31__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_38__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_45__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_52__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_59__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_66__pin_a2f_o_0_, chanx_right_in[83]}),
		.sram(mux_tree_tapbuf_L4SB_size8_54_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_54_sram_inv[0:2]),
		.out(chany_top_out[82]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_166 (
		.in({top_right_grid_left_width_0_height_0_subtile_25__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_32__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_39__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_46__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_53__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_60__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_67__pin_a2f_o_0_, chanx_right_in[84]}),
		.sram(mux_tree_tapbuf_L4SB_size8_55_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_55_sram_inv[0:2]),
		.out(chany_top_out[83]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_168 (
		.in({top_right_grid_left_width_0_height_0_subtile_26__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_33__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_40__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_47__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_54__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_61__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_68__pin_a2f_o_0_, chanx_right_in[85]}),
		.sram(mux_tree_tapbuf_L4SB_size8_56_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_56_sram_inv[0:2]),
		.out(chany_top_out[84]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_170 (
		.in({top_right_grid_left_width_0_height_0_subtile_27__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_34__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_41__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_48__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_55__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_62__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_69__pin_a2f_o_0_, chanx_right_in[86]}),
		.sram(mux_tree_tapbuf_L4SB_size8_57_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_57_sram_inv[0:2]),
		.out(chany_top_out[85]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_172 (
		.in({top_right_grid_left_width_0_height_0_subtile_28__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_35__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_42__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_49__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_56__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_63__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_70__pin_a2f_o_0_, chanx_right_in[87]}),
		.sram(mux_tree_tapbuf_L4SB_size8_58_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_58_sram_inv[0:2]),
		.out(chany_top_out[86]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_174 (
		.in({top_right_grid_left_width_0_height_0_subtile_29__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_36__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_43__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_50__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_57__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_64__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_71__pin_a2f_o_0_, chanx_right_in[88]}),
		.sram(mux_tree_tapbuf_L4SB_size8_59_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_59_sram_inv[0:2]),
		.out(chany_top_out[87]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_178 (
		.in({top_right_grid_left_width_0_height_0_subtile_24__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_31__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_38__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_45__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_52__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_59__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_66__pin_a2f_o_0_, chanx_right_in[90]}),
		.sram(mux_tree_tapbuf_L4SB_size8_60_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_60_sram_inv[0:2]),
		.out(chany_top_out[89]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_180 (
		.in({top_right_grid_left_width_0_height_0_subtile_25__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_32__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_39__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_46__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_53__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_60__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_67__pin_a2f_o_0_, chanx_right_in[91]}),
		.sram(mux_tree_tapbuf_L4SB_size8_61_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_61_sram_inv[0:2]),
		.out(chany_top_out[90]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_182 (
		.in({top_right_grid_left_width_0_height_0_subtile_26__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_33__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_40__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_47__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_54__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_61__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_68__pin_a2f_o_0_, chanx_right_in[92]}),
		.sram(mux_tree_tapbuf_L4SB_size8_62_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_62_sram_inv[0:2]),
		.out(chany_top_out[91]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_184 (
		.in({top_right_grid_left_width_0_height_0_subtile_27__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_34__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_41__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_48__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_55__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_62__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_69__pin_a2f_o_0_, chanx_right_in[93]}),
		.sram(mux_tree_tapbuf_L4SB_size8_63_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_63_sram_inv[0:2]),
		.out(chany_top_out[92]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_186 (
		.in({top_right_grid_left_width_0_height_0_subtile_28__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_35__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_42__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_49__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_56__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_63__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_70__pin_a2f_o_0_, chanx_right_in[94]}),
		.sram(mux_tree_tapbuf_L4SB_size8_64_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_64_sram_inv[0:2]),
		.out(chany_top_out[93]));

	mux_tree_tapbuf_L4SB_size8 mux_top_track_188 (
		.in({top_right_grid_left_width_0_height_0_subtile_29__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_36__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_43__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_50__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_57__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_64__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_71__pin_a2f_o_0_, chanx_right_in[95]}),
		.sram(mux_tree_tapbuf_L4SB_size8_65_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_65_sram_inv[0:2]),
		.out(chany_top_out[94]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_38 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size3_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_0_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_40 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_1_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_42 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_2_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_44 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_3_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_46 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_4_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_4_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_48 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_5_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_5_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_52 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size7_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_6_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_6_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_54 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_7_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_7_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_56 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_8_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_8_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_58 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_9_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_9_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_60 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_10_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_10_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_62 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_11_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_11_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_66 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size7_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_12_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_12_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_68 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_13_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_13_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_70 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_14_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_14_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_72 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_15_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_15_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_74 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_16_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_16_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_76 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_17_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_17_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_80 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size7_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_18_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_18_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_82 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_19_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_19_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_84 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_20_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_20_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_86 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_21_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_21_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_88 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_22_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_22_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_90 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_23_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_23_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_94 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size7_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_24_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_24_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_96 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_25_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_25_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_98 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_26_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_26_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_100 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_27_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_27_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_27_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_102 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_27_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_28_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_28_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_28_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_104 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_28_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_29_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_29_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_29_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_108 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size7_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_30_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_30_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_30_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_110 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_30_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_31_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_31_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_31_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_112 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_31_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_32_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_32_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_32_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_114 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_32_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_33_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_33_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_33_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_116 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_33_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_34_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_34_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_34_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_118 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_34_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_35_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_35_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_35_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_122 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size7_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_36_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_36_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_36_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_124 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_36_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_37_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_37_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_37_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_126 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_37_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_38_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_38_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_38_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_128 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_38_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_39_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_39_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_39_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_130 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_39_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_40_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_40_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_40_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_132 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_40_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_41_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_41_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_41_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_136 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size7_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_42_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_42_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_42_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_138 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_42_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_43_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_43_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_43_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_140 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_43_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_44_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_44_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_44_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_142 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_44_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_45_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_45_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_45_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_144 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_45_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_46_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_46_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_46_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_146 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_46_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_47_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_47_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_47_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_150 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size7_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_48_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_48_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_48_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_152 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_48_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_49_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_49_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_49_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_154 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_49_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_50_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_50_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_50_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_156 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_50_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_51_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_51_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_51_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_158 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_51_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_52_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_52_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_52_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_160 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_52_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_53_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_53_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_53_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_164 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size7_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_54_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_54_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_54_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_166 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_54_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_55_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_55_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_55_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_168 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_55_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_56_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_56_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_56_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_170 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_56_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_57_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_57_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_57_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_172 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_57_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_58_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_58_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_58_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_174 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_58_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_59_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_59_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_59_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_178 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size7_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_60_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_60_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_60_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_180 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_60_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_61_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_61_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_61_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_182 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_61_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_62_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_62_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_62_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_184 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_62_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_63_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_63_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_63_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_186 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_63_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_64_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_64_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_64_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_top_track_188 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_64_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_65_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_65_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_65_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7 mux_top_track_50 (
		.in({top_right_grid_left_width_0_height_0_subtile_30__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_37__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_44__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_51__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_58__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_65__pin_a2f_o_0_, chanx_right_in[26]}),
		.sram(mux_tree_tapbuf_L4SB_size7_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_0_sram_inv[0:2]),
		.out(chany_top_out[25]));

	mux_tree_tapbuf_L4SB_size7 mux_top_track_64 (
		.in({top_right_grid_left_width_0_height_0_subtile_30__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_37__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_44__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_51__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_58__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_65__pin_a2f_o_0_, chanx_right_in[33]}),
		.sram(mux_tree_tapbuf_L4SB_size7_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_1_sram_inv[0:2]),
		.out(chany_top_out[32]));

	mux_tree_tapbuf_L4SB_size7 mux_top_track_78 (
		.in({top_right_grid_left_width_0_height_0_subtile_30__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_37__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_44__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_51__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_58__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_65__pin_a2f_o_0_, chanx_right_in[40]}),
		.sram(mux_tree_tapbuf_L4SB_size7_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_2_sram_inv[0:2]),
		.out(chany_top_out[39]));

	mux_tree_tapbuf_L4SB_size7 mux_top_track_92 (
		.in({top_right_grid_left_width_0_height_0_subtile_30__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_37__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_44__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_51__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_58__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_65__pin_a2f_o_0_, chanx_right_in[47]}),
		.sram(mux_tree_tapbuf_L4SB_size7_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_3_sram_inv[0:2]),
		.out(chany_top_out[46]));

	mux_tree_tapbuf_L4SB_size7 mux_top_track_106 (
		.in({top_right_grid_left_width_0_height_0_subtile_30__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_37__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_44__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_51__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_58__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_65__pin_a2f_o_0_, chanx_right_in[54]}),
		.sram(mux_tree_tapbuf_L4SB_size7_4_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_4_sram_inv[0:2]),
		.out(chany_top_out[53]));

	mux_tree_tapbuf_L4SB_size7 mux_top_track_120 (
		.in({top_right_grid_left_width_0_height_0_subtile_30__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_37__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_44__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_51__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_58__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_65__pin_a2f_o_0_, chanx_right_in[61]}),
		.sram(mux_tree_tapbuf_L4SB_size7_5_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_5_sram_inv[0:2]),
		.out(chany_top_out[60]));

	mux_tree_tapbuf_L4SB_size7 mux_top_track_134 (
		.in({top_right_grid_left_width_0_height_0_subtile_30__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_37__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_44__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_51__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_58__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_65__pin_a2f_o_0_, chanx_right_in[68]}),
		.sram(mux_tree_tapbuf_L4SB_size7_6_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_6_sram_inv[0:2]),
		.out(chany_top_out[67]));

	mux_tree_tapbuf_L4SB_size7 mux_top_track_148 (
		.in({top_right_grid_left_width_0_height_0_subtile_30__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_37__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_44__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_51__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_58__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_65__pin_a2f_o_0_, chanx_right_in[75]}),
		.sram(mux_tree_tapbuf_L4SB_size7_7_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_7_sram_inv[0:2]),
		.out(chany_top_out[74]));

	mux_tree_tapbuf_L4SB_size7 mux_top_track_162 (
		.in({top_right_grid_left_width_0_height_0_subtile_30__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_37__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_44__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_51__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_58__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_65__pin_a2f_o_0_, chanx_right_in[82]}),
		.sram(mux_tree_tapbuf_L4SB_size7_8_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_8_sram_inv[0:2]),
		.out(chany_top_out[81]));

	mux_tree_tapbuf_L4SB_size7 mux_top_track_176 (
		.in({top_right_grid_left_width_0_height_0_subtile_30__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_37__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_44__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_51__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_58__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_65__pin_a2f_o_0_, chanx_right_in[89]}),
		.sram(mux_tree_tapbuf_L4SB_size7_9_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_9_sram_inv[0:2]),
		.out(chany_top_out[88]));

	mux_tree_tapbuf_L4SB_size7 mux_top_track_190 (
		.in({top_right_grid_left_width_0_height_0_subtile_30__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_37__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_44__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_51__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_58__pin_a2f_o_0_, top_right_grid_left_width_0_height_0_subtile_65__pin_a2f_o_0_, chanx_right_in[0]}),
		.sram(mux_tree_tapbuf_L4SB_size7_10_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_10_sram_inv[0:2]),
		.out(chany_top_out[95]));

	mux_tree_tapbuf_L4SB_size7_mem mem_top_track_50 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size7_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size7_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_0_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7_mem mem_top_track_64 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size7_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size7_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_1_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7_mem mem_top_track_78 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size7_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size7_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_2_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7_mem mem_top_track_92 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size7_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size7_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_3_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7_mem mem_top_track_106 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_29_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size7_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size7_4_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_4_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7_mem mem_top_track_120 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_35_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size7_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size7_5_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_5_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7_mem mem_top_track_134 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_41_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size7_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size7_6_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_6_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7_mem mem_top_track_148 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_47_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size7_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size7_7_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_7_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7_mem mem_top_track_162 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_53_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size7_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size7_8_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_8_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7_mem mem_top_track_176 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_59_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size7_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size7_9_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_9_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7_mem mem_top_track_190 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_65_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size7_10_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_10_sram_inv[0:2]));

endmodule
// ----- END Verilog module for sb_0__0_ -----

//----- Default net type -----
`default_nettype none



