//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for Unique Switch Blocks[10][8]
//	Author: Xifan TANG
//	Organization: University of Utah
//-------------------------------------------
//----- Time scale -----
`timescale 1ns / 1ps

//----- Default net type -----
`default_nettype wire

// ----- Verilog module for sb_10__8_ -----
module sb_10__8_(config_enable,
                 prog_clock,
                 chany_bottom_in,
                 bottom_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_1_,
                 bottom_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_1_,
                 bottom_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_1_,
                 bottom_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_1_,
                 bottom_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_1_,
                 bottom_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_1_,
                 bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_1_,
                 bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_1_,
                 bottom_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_1_,
                 bottom_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_1_,
                 bottom_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_1_,
                 bottom_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_1_,
                 bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_1_,
                 bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_1_,
                 bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_1_,
                 bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_1_,
                 bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_1_,
                 bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_1_,
                 bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_1_,
                 bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_1_,
                 bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_1_,
                 bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_1_,
                 bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_1_,
                 bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_1_,
                 bottom_left_grid_right_width_0_height_0_subtile_24__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_24__pin_a2f_o_1_,
                 bottom_left_grid_right_width_0_height_0_subtile_25__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_25__pin_a2f_o_1_,
                 bottom_left_grid_right_width_0_height_0_subtile_26__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_26__pin_a2f_o_1_,
                 bottom_left_grid_right_width_0_height_0_subtile_27__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_27__pin_a2f_o_1_,
                 bottom_left_grid_right_width_0_height_0_subtile_28__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_28__pin_a2f_o_1_,
                 bottom_left_grid_right_width_0_height_0_subtile_29__pin_a2f_o_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_29__pin_a2f_o_1_,
                 chanx_left_in,
                 left_bottom_grid_top_width_0_height_0_subtile_30__pin_a2f_o_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_30__pin_a2f_o_1_,
                 left_bottom_grid_top_width_0_height_0_subtile_31__pin_a2f_o_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_31__pin_a2f_o_1_,
                 left_bottom_grid_top_width_0_height_0_subtile_32__pin_a2f_o_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_32__pin_a2f_o_1_,
                 left_bottom_grid_top_width_0_height_0_subtile_33__pin_a2f_o_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_33__pin_a2f_o_1_,
                 left_bottom_grid_top_width_0_height_0_subtile_34__pin_a2f_o_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_34__pin_a2f_o_1_,
                 left_bottom_grid_top_width_0_height_0_subtile_35__pin_a2f_o_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_35__pin_a2f_o_1_,
                 left_bottom_grid_top_width_0_height_0_subtile_36__pin_a2f_o_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_36__pin_a2f_o_1_,
                 left_bottom_grid_top_width_0_height_0_subtile_37__pin_a2f_o_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_37__pin_a2f_o_1_,
                 left_bottom_grid_top_width_0_height_0_subtile_38__pin_a2f_o_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_38__pin_a2f_o_1_,
                 left_bottom_grid_top_width_0_height_0_subtile_39__pin_a2f_o_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_39__pin_a2f_o_1_,
                 left_bottom_grid_top_width_0_height_0_subtile_40__pin_a2f_o_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_40__pin_a2f_o_1_,
                 left_bottom_grid_top_width_0_height_0_subtile_41__pin_a2f_o_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_41__pin_a2f_o_1_,
                 left_bottom_grid_top_width_0_height_0_subtile_42__pin_a2f_o_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_42__pin_a2f_o_1_,
                 left_bottom_grid_top_width_0_height_0_subtile_43__pin_a2f_o_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_43__pin_a2f_o_1_,
                 left_bottom_grid_top_width_0_height_0_subtile_44__pin_a2f_o_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_44__pin_a2f_o_1_,
                 left_bottom_grid_top_width_0_height_0_subtile_45__pin_a2f_o_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_45__pin_a2f_o_1_,
                 left_bottom_grid_top_width_0_height_0_subtile_46__pin_a2f_o_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_46__pin_a2f_o_1_,
                 left_bottom_grid_top_width_0_height_0_subtile_47__pin_a2f_o_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_47__pin_a2f_o_1_,
                 left_bottom_grid_top_width_0_height_0_subtile_48__pin_a2f_o_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_48__pin_a2f_o_1_,
                 left_bottom_grid_top_width_0_height_0_subtile_49__pin_a2f_o_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_49__pin_a2f_o_1_,
                 left_bottom_grid_top_width_0_height_0_subtile_50__pin_a2f_o_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_50__pin_a2f_o_1_,
                 left_bottom_grid_top_width_0_height_0_subtile_51__pin_a2f_o_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_51__pin_a2f_o_1_,
                 left_bottom_grid_top_width_0_height_0_subtile_52__pin_a2f_o_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_52__pin_a2f_o_1_,
                 left_bottom_grid_top_width_0_height_0_subtile_53__pin_a2f_o_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_53__pin_a2f_o_1_,
                 left_bottom_grid_top_width_0_height_0_subtile_54__pin_a2f_o_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_54__pin_a2f_o_1_,
                 left_bottom_grid_top_width_0_height_0_subtile_55__pin_a2f_o_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_55__pin_a2f_o_1_,
                 left_bottom_grid_top_width_0_height_0_subtile_56__pin_a2f_o_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_56__pin_a2f_o_1_,
                 left_bottom_grid_top_width_0_height_0_subtile_57__pin_a2f_o_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_57__pin_a2f_o_1_,
                 left_bottom_grid_top_width_0_height_0_subtile_58__pin_a2f_o_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_58__pin_a2f_o_1_,
                 left_bottom_grid_top_width_0_height_0_subtile_59__pin_a2f_o_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_59__pin_a2f_o_1_,
                 ccff_head,
                 chany_bottom_out,
                 chanx_left_out,
                 ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_clock;
//----- INPUT PORTS -----
input [0:95] chany_bottom_in;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_24__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_24__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_25__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_25__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_26__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_26__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_27__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_27__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_28__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_28__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_29__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_29__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:95] chanx_left_in;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_30__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_30__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_31__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_31__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_32__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_32__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_33__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_33__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_34__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_34__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_35__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_35__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_36__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_36__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_37__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_37__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_38__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_38__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_39__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_39__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_40__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_40__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_41__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_41__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_42__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_42__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_43__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_43__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_44__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_44__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_45__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_45__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_46__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_46__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_47__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_47__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_48__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_48__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_49__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_49__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_50__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_50__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_51__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_51__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_52__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_52__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_53__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_53__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_54__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_54__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_55__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_55__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_56__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_56__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_57__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_57__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_58__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_58__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_59__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_59__pin_a2f_o_1_;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:95] chany_bottom_out;
//----- OUTPUT PORTS -----
output [0:95] chanx_left_out;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:1] mux_tree_tapbuf_L2SB_size4_0_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_0_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_10_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_10_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_11_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_11_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_12_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_12_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_13_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_13_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_14_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_14_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_15_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_15_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_16_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_16_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_17_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_17_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_18_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_18_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_19_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_19_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_1_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_1_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_20_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_20_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_21_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_21_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_22_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_22_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_23_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_23_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_24_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_24_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_25_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_25_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_26_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_26_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_27_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_27_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_28_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_28_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_29_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_29_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_2_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_2_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_30_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_30_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_31_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_31_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_3_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_3_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_4_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_4_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_5_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_5_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_6_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_6_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_7_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_7_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_8_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_8_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_9_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_9_sram_inv;
wire [0:2] mux_tree_tapbuf_L2SB_size5_0_sram;
wire [0:2] mux_tree_tapbuf_L2SB_size5_0_sram_inv;
wire [0:2] mux_tree_tapbuf_L2SB_size5_1_sram;
wire [0:2] mux_tree_tapbuf_L2SB_size5_1_sram_inv;
wire [0:2] mux_tree_tapbuf_L2SB_size5_2_sram;
wire [0:2] mux_tree_tapbuf_L2SB_size5_2_sram_inv;
wire [0:2] mux_tree_tapbuf_L2SB_size5_3_sram;
wire [0:2] mux_tree_tapbuf_L2SB_size5_3_sram_inv;
wire [0:2] mux_tree_tapbuf_L2SB_size5_4_sram;
wire [0:2] mux_tree_tapbuf_L2SB_size5_4_sram_inv;
wire [0:2] mux_tree_tapbuf_L2SB_size5_5_sram;
wire [0:2] mux_tree_tapbuf_L2SB_size5_5_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size10_0_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size10_0_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size10_10_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size10_10_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size10_11_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size10_11_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size10_12_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size10_12_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size10_13_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size10_13_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size10_1_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size10_1_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size10_2_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size10_2_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size10_3_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size10_3_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size10_4_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size10_4_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size10_5_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size10_5_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size10_6_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size10_6_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size10_7_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size10_7_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size10_8_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size10_8_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size10_9_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size10_9_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size11_0_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size11_0_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size11_10_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size11_10_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size11_11_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size11_11_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size11_12_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size11_12_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size11_13_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size11_13_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size11_14_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size11_14_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size11_15_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size11_15_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size11_16_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size11_16_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size11_17_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size11_17_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size11_18_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size11_18_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size11_19_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size11_19_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size11_1_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size11_1_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size11_2_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size11_2_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size11_3_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size11_3_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size11_4_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size11_4_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size11_5_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size11_5_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size11_6_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size11_6_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size11_7_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size11_7_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size11_8_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size11_8_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size11_9_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size11_9_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size12_0_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size12_0_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size12_10_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size12_10_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size12_11_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size12_11_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size12_12_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size12_12_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size12_13_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size12_13_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size12_14_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size12_14_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size12_15_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size12_15_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size12_1_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size12_1_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size12_2_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size12_2_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size12_3_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size12_3_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size12_4_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size12_4_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size12_5_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size12_5_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size12_6_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size12_6_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size12_7_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size12_7_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size12_8_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size12_8_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size12_9_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size12_9_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size13_0_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size13_0_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size13_10_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size13_10_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size13_11_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size13_11_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size13_12_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size13_12_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size13_13_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size13_13_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size13_14_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size13_14_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size13_15_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size13_15_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size13_16_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size13_16_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size13_17_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size13_17_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size13_18_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size13_18_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size13_19_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size13_19_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size13_1_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size13_1_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size13_2_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size13_2_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size13_3_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size13_3_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size13_4_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size13_4_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size13_5_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size13_5_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size13_6_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size13_6_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size13_7_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size13_7_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size13_8_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size13_8_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size13_9_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size13_9_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size14_0_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size14_0_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size14_1_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size14_1_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_0_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_0_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_10_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_10_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_11_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_11_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_12_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_12_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_13_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_13_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_1_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_1_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_2_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_2_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_3_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_3_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_4_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_4_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_5_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_5_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_6_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_6_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_7_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_7_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_8_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_8_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size5_9_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size5_9_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size6_0_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size6_0_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size6_10_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size6_10_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size6_11_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size6_11_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size6_12_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size6_12_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size6_13_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size6_13_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size6_14_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size6_14_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size6_15_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size6_15_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size6_16_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size6_16_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size6_17_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size6_17_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size6_18_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size6_18_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size6_19_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size6_19_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size6_1_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size6_1_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size6_20_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size6_20_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size6_21_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size6_21_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size6_2_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size6_2_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size6_3_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size6_3_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size6_4_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size6_4_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size6_5_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size6_5_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size6_6_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size6_6_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size6_7_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size6_7_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size6_8_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size6_8_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size6_9_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size6_9_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_0_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_0_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_10_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_10_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_11_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_11_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_1_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_1_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_2_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_2_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_3_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_3_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_4_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_4_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_5_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_5_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_6_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_6_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_7_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_7_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_8_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_8_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_9_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_9_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_0_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_0_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_10_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_10_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_11_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_11_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_12_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_12_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_13_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_13_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_14_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_14_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_15_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_15_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_16_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_16_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_17_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_17_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_1_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_1_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_2_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_2_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_3_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_3_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_4_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_4_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_5_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_5_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_6_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_6_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_7_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_7_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_8_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_8_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_9_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_9_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_0_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_0_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_10_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_10_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_11_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_11_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_12_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_12_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_13_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_13_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_14_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_14_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_15_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_15_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_1_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_1_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_2_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_2_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_3_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_3_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_4_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_4_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_5_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_5_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_6_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_6_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_7_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_7_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_8_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_8_sram_inv;
wire [0:3] mux_tree_tapbuf_L4SB_size9_9_sram;
wire [0:3] mux_tree_tapbuf_L4SB_size9_9_sram_inv;

// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	mux_tree_tapbuf_L2SB_size5 mux_bottom_track_1 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_28__pin_a2f_o_1_, chanx_left_in[1]}),
		.sram(mux_tree_tapbuf_L2SB_size5_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L2SB_size5_0_sram_inv[0:2]),
		.out(chany_bottom_out[0]));

	mux_tree_tapbuf_L2SB_size5 mux_bottom_track_3 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_29__pin_a2f_o_0_, chanx_left_in[2]}),
		.sram(mux_tree_tapbuf_L2SB_size5_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L2SB_size5_1_sram_inv[0:2]),
		.out(chany_bottom_out[1]));

	mux_tree_tapbuf_L2SB_size5 mux_bottom_track_5 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_29__pin_a2f_o_1_, chanx_left_in[3]}),
		.sram(mux_tree_tapbuf_L2SB_size5_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L2SB_size5_2_sram_inv[0:2]),
		.out(chany_bottom_out[2]));

	mux_tree_tapbuf_L2SB_size5 mux_left_track_1 (
		.in({chany_bottom_in[95], left_bottom_grid_top_width_0_height_0_subtile_30__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_39__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_49__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_58__pin_a2f_o_1_}),
		.sram(mux_tree_tapbuf_L2SB_size5_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L2SB_size5_3_sram_inv[0:2]),
		.out(chanx_left_out[0]));

	mux_tree_tapbuf_L2SB_size5 mux_left_track_3 (
		.in({chany_bottom_in[0], left_bottom_grid_top_width_0_height_0_subtile_30__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_40__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_49__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_59__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L2SB_size5_4_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L2SB_size5_4_sram_inv[0:2]),
		.out(chanx_left_out[1]));

	mux_tree_tapbuf_L2SB_size5 mux_left_track_5 (
		.in({chany_bottom_in[1], left_bottom_grid_top_width_0_height_0_subtile_31__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_40__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_50__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_59__pin_a2f_o_1_}),
		.sram(mux_tree_tapbuf_L2SB_size5_5_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L2SB_size5_5_sram_inv[0:2]),
		.out(chanx_left_out[2]));

	mux_tree_tapbuf_L2SB_size5_mem mem_bottom_track_1 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(ccff_head),
		.ccff_tail(mux_tree_tapbuf_L2SB_size5_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size5_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L2SB_size5_0_sram_inv[0:2]));

	mux_tree_tapbuf_L2SB_size5_mem mem_bottom_track_3 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size5_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size5_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size5_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L2SB_size5_1_sram_inv[0:2]));

	mux_tree_tapbuf_L2SB_size5_mem mem_bottom_track_5 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size5_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size5_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size5_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L2SB_size5_2_sram_inv[0:2]));

	mux_tree_tapbuf_L2SB_size5_mem mem_left_track_1 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size5_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size5_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size5_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L2SB_size5_3_sram_inv[0:2]));

	mux_tree_tapbuf_L2SB_size5_mem mem_left_track_3 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size5_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size5_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size5_4_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L2SB_size5_4_sram_inv[0:2]));

	mux_tree_tapbuf_L2SB_size5_mem mem_left_track_5 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size5_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size5_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size5_5_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L2SB_size5_5_sram_inv[0:2]));

	mux_tree_tapbuf_L2SB_size4 mux_bottom_track_7 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_1_, chanx_left_in[4]}),
		.sram(mux_tree_tapbuf_L2SB_size4_0_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_0_sram_inv[0:1]),
		.out(chany_bottom_out[3]));

	mux_tree_tapbuf_L2SB_size4 mux_bottom_track_9 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_, chanx_left_in[5]}),
		.sram(mux_tree_tapbuf_L2SB_size4_1_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_1_sram_inv[0:1]),
		.out(chany_bottom_out[4]));

	mux_tree_tapbuf_L2SB_size4 mux_bottom_track_11 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_1_, chanx_left_in[6]}),
		.sram(mux_tree_tapbuf_L2SB_size4_2_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_2_sram_inv[0:1]),
		.out(chany_bottom_out[5]));

	mux_tree_tapbuf_L2SB_size4 mux_bottom_track_13 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_, chanx_left_in[7]}),
		.sram(mux_tree_tapbuf_L2SB_size4_3_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_3_sram_inv[0:1]),
		.out(chany_bottom_out[6]));

	mux_tree_tapbuf_L2SB_size4 mux_bottom_track_15 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_1_, chanx_left_in[8]}),
		.sram(mux_tree_tapbuf_L2SB_size4_4_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_4_sram_inv[0:1]),
		.out(chany_bottom_out[7]));

	mux_tree_tapbuf_L2SB_size4 mux_bottom_track_17 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_, chanx_left_in[9]}),
		.sram(mux_tree_tapbuf_L2SB_size4_5_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_5_sram_inv[0:1]),
		.out(chany_bottom_out[8]));

	mux_tree_tapbuf_L2SB_size4 mux_bottom_track_19 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_1_, chanx_left_in[10]}),
		.sram(mux_tree_tapbuf_L2SB_size4_6_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_6_sram_inv[0:1]),
		.out(chany_bottom_out[9]));

	mux_tree_tapbuf_L2SB_size4 mux_bottom_track_21 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_24__pin_a2f_o_0_, chanx_left_in[11]}),
		.sram(mux_tree_tapbuf_L2SB_size4_7_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_7_sram_inv[0:1]),
		.out(chany_bottom_out[10]));

	mux_tree_tapbuf_L2SB_size4 mux_bottom_track_23 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_24__pin_a2f_o_1_, chanx_left_in[12]}),
		.sram(mux_tree_tapbuf_L2SB_size4_8_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_8_sram_inv[0:1]),
		.out(chany_bottom_out[11]));

	mux_tree_tapbuf_L2SB_size4 mux_bottom_track_25 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_25__pin_a2f_o_0_, chanx_left_in[13]}),
		.sram(mux_tree_tapbuf_L2SB_size4_9_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_9_sram_inv[0:1]),
		.out(chany_bottom_out[12]));

	mux_tree_tapbuf_L2SB_size4 mux_bottom_track_27 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_25__pin_a2f_o_1_, chanx_left_in[14]}),
		.sram(mux_tree_tapbuf_L2SB_size4_10_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_10_sram_inv[0:1]),
		.out(chany_bottom_out[13]));

	mux_tree_tapbuf_L2SB_size4 mux_bottom_track_29 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_26__pin_a2f_o_0_, chanx_left_in[15]}),
		.sram(mux_tree_tapbuf_L2SB_size4_11_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_11_sram_inv[0:1]),
		.out(chany_bottom_out[14]));

	mux_tree_tapbuf_L2SB_size4 mux_bottom_track_31 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_26__pin_a2f_o_1_, chanx_left_in[16]}),
		.sram(mux_tree_tapbuf_L2SB_size4_12_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_12_sram_inv[0:1]),
		.out(chany_bottom_out[15]));

	mux_tree_tapbuf_L2SB_size4 mux_bottom_track_33 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_27__pin_a2f_o_0_, chanx_left_in[17]}),
		.sram(mux_tree_tapbuf_L2SB_size4_13_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_13_sram_inv[0:1]),
		.out(chany_bottom_out[16]));

	mux_tree_tapbuf_L2SB_size4 mux_bottom_track_35 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_27__pin_a2f_o_1_, chanx_left_in[18]}),
		.sram(mux_tree_tapbuf_L2SB_size4_14_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_14_sram_inv[0:1]),
		.out(chany_bottom_out[17]));

	mux_tree_tapbuf_L2SB_size4 mux_bottom_track_37 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_28__pin_a2f_o_0_, chanx_left_in[19]}),
		.sram(mux_tree_tapbuf_L2SB_size4_15_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_15_sram_inv[0:1]),
		.out(chany_bottom_out[18]));

	mux_tree_tapbuf_L2SB_size4 mux_left_track_7 (
		.in({chany_bottom_in[2], left_bottom_grid_top_width_0_height_0_subtile_31__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_41__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_50__pin_a2f_o_1_}),
		.sram(mux_tree_tapbuf_L2SB_size4_16_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_16_sram_inv[0:1]),
		.out(chanx_left_out[3]));

	mux_tree_tapbuf_L2SB_size4 mux_left_track_9 (
		.in({chany_bottom_in[3], left_bottom_grid_top_width_0_height_0_subtile_32__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_41__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_51__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L2SB_size4_17_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_17_sram_inv[0:1]),
		.out(chanx_left_out[4]));

	mux_tree_tapbuf_L2SB_size4 mux_left_track_11 (
		.in({chany_bottom_in[4], left_bottom_grid_top_width_0_height_0_subtile_32__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_42__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_51__pin_a2f_o_1_}),
		.sram(mux_tree_tapbuf_L2SB_size4_18_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_18_sram_inv[0:1]),
		.out(chanx_left_out[5]));

	mux_tree_tapbuf_L2SB_size4 mux_left_track_13 (
		.in({chany_bottom_in[5], left_bottom_grid_top_width_0_height_0_subtile_33__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_42__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_52__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L2SB_size4_19_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_19_sram_inv[0:1]),
		.out(chanx_left_out[6]));

	mux_tree_tapbuf_L2SB_size4 mux_left_track_15 (
		.in({chany_bottom_in[6], left_bottom_grid_top_width_0_height_0_subtile_33__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_43__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_52__pin_a2f_o_1_}),
		.sram(mux_tree_tapbuf_L2SB_size4_20_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_20_sram_inv[0:1]),
		.out(chanx_left_out[7]));

	mux_tree_tapbuf_L2SB_size4 mux_left_track_17 (
		.in({chany_bottom_in[7], left_bottom_grid_top_width_0_height_0_subtile_34__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_43__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_53__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L2SB_size4_21_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_21_sram_inv[0:1]),
		.out(chanx_left_out[8]));

	mux_tree_tapbuf_L2SB_size4 mux_left_track_19 (
		.in({chany_bottom_in[8], left_bottom_grid_top_width_0_height_0_subtile_34__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_44__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_53__pin_a2f_o_1_}),
		.sram(mux_tree_tapbuf_L2SB_size4_22_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_22_sram_inv[0:1]),
		.out(chanx_left_out[9]));

	mux_tree_tapbuf_L2SB_size4 mux_left_track_21 (
		.in({chany_bottom_in[9], left_bottom_grid_top_width_0_height_0_subtile_35__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_44__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_54__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L2SB_size4_23_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_23_sram_inv[0:1]),
		.out(chanx_left_out[10]));

	mux_tree_tapbuf_L2SB_size4 mux_left_track_23 (
		.in({chany_bottom_in[10], left_bottom_grid_top_width_0_height_0_subtile_35__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_45__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_54__pin_a2f_o_1_}),
		.sram(mux_tree_tapbuf_L2SB_size4_24_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_24_sram_inv[0:1]),
		.out(chanx_left_out[11]));

	mux_tree_tapbuf_L2SB_size4 mux_left_track_25 (
		.in({chany_bottom_in[11], left_bottom_grid_top_width_0_height_0_subtile_36__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_45__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_55__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L2SB_size4_25_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_25_sram_inv[0:1]),
		.out(chanx_left_out[12]));

	mux_tree_tapbuf_L2SB_size4 mux_left_track_27 (
		.in({chany_bottom_in[12], left_bottom_grid_top_width_0_height_0_subtile_36__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_46__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_55__pin_a2f_o_1_}),
		.sram(mux_tree_tapbuf_L2SB_size4_26_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_26_sram_inv[0:1]),
		.out(chanx_left_out[13]));

	mux_tree_tapbuf_L2SB_size4 mux_left_track_29 (
		.in({chany_bottom_in[13], left_bottom_grid_top_width_0_height_0_subtile_37__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_46__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_56__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L2SB_size4_27_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_27_sram_inv[0:1]),
		.out(chanx_left_out[14]));

	mux_tree_tapbuf_L2SB_size4 mux_left_track_31 (
		.in({chany_bottom_in[14], left_bottom_grid_top_width_0_height_0_subtile_37__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_47__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_56__pin_a2f_o_1_}),
		.sram(mux_tree_tapbuf_L2SB_size4_28_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_28_sram_inv[0:1]),
		.out(chanx_left_out[15]));

	mux_tree_tapbuf_L2SB_size4 mux_left_track_33 (
		.in({chany_bottom_in[15], left_bottom_grid_top_width_0_height_0_subtile_38__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_47__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_57__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L2SB_size4_29_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_29_sram_inv[0:1]),
		.out(chanx_left_out[16]));

	mux_tree_tapbuf_L2SB_size4 mux_left_track_35 (
		.in({chany_bottom_in[16], left_bottom_grid_top_width_0_height_0_subtile_38__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_48__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_57__pin_a2f_o_1_}),
		.sram(mux_tree_tapbuf_L2SB_size4_30_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_30_sram_inv[0:1]),
		.out(chanx_left_out[17]));

	mux_tree_tapbuf_L2SB_size4 mux_left_track_37 (
		.in({chany_bottom_in[17], left_bottom_grid_top_width_0_height_0_subtile_39__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_48__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_58__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L2SB_size4_31_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_31_sram_inv[0:1]),
		.out(chanx_left_out[18]));

	mux_tree_tapbuf_L2SB_size4_mem mem_bottom_track_7 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size5_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_0_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_0_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_bottom_track_9 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_1_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_1_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_bottom_track_11 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_2_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_2_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_bottom_track_13 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_3_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_3_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_bottom_track_15 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_4_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_4_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_bottom_track_17 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_5_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_5_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_bottom_track_19 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_6_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_6_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_bottom_track_21 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_7_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_7_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_bottom_track_23 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_8_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_8_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_bottom_track_25 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_9_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_9_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_bottom_track_27 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_10_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_10_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_bottom_track_29 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_11_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_11_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_bottom_track_31 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_12_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_12_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_bottom_track_33 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_13_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_13_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_bottom_track_35 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_14_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_14_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_bottom_track_37 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_15_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_15_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_left_track_7 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size5_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_16_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_16_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_left_track_9 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_17_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_17_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_left_track_11 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_18_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_18_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_left_track_13 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_19_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_19_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_left_track_15 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_20_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_20_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_left_track_17 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_21_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_21_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_left_track_19 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_22_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_22_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_left_track_21 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_23_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_23_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_left_track_23 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_24_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_24_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_left_track_25 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_25_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_25_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_left_track_27 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_26_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_26_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_left_track_29 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_27_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_27_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_27_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_left_track_31 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_27_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_28_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_28_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_28_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_left_track_33 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_28_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_29_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_29_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_29_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_left_track_35 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_29_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_30_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_30_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_30_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_left_track_37 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_30_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_31_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_31_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_31_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size13 mux_bottom_track_39 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_26__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_28__pin_a2f_o_0_, chanx_left_in[20]}),
		.sram(mux_tree_tapbuf_L4SB_size13_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size13_0_sram_inv[0:3]),
		.out(chany_bottom_out[19]));

	mux_tree_tapbuf_L4SB_size13 mux_bottom_track_43 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_27__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_29__pin_a2f_o_0_, chanx_left_in[22]}),
		.sram(mux_tree_tapbuf_L4SB_size13_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size13_1_sram_inv[0:3]),
		.out(chany_bottom_out[21]));

	mux_tree_tapbuf_L4SB_size13 mux_bottom_track_137 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_24__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_28__pin_a2f_o_0_, chanx_left_in[69]}),
		.sram(mux_tree_tapbuf_L4SB_size13_2_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size13_2_sram_inv[0:3]),
		.out(chany_bottom_out[68]));

	mux_tree_tapbuf_L4SB_size13 mux_bottom_track_141 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_25__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_29__pin_a2f_o_0_, chanx_left_in[71]}),
		.sram(mux_tree_tapbuf_L4SB_size13_3_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size13_3_sram_inv[0:3]),
		.out(chany_bottom_out[70]));

	mux_tree_tapbuf_L4SB_size13 mux_bottom_track_153 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_24__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_25__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_28__pin_a2f_o_1_, chanx_left_in[77]}),
		.sram(mux_tree_tapbuf_L4SB_size13_4_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size13_4_sram_inv[0:3]),
		.out(chany_bottom_out[76]));

	mux_tree_tapbuf_L4SB_size13 mux_bottom_track_157 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_25__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_26__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_29__pin_a2f_o_1_, chanx_left_in[79]}),
		.sram(mux_tree_tapbuf_L4SB_size13_5_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size13_5_sram_inv[0:3]),
		.out(chany_bottom_out[78]));

	mux_tree_tapbuf_L4SB_size13 mux_bottom_track_165 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_27__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_28__pin_a2f_o_0_, chanx_left_in[83]}),
		.sram(mux_tree_tapbuf_L4SB_size13_6_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size13_6_sram_inv[0:3]),
		.out(chany_bottom_out[82]));

	mux_tree_tapbuf_L4SB_size13 mux_bottom_track_173 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_25__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_29__pin_a2f_o_1_, chanx_left_in[87]}),
		.sram(mux_tree_tapbuf_L4SB_size13_7_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size13_7_sram_inv[0:3]),
		.out(chany_bottom_out[86]));

	mux_tree_tapbuf_L4SB_size13 mux_bottom_track_185 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_24__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_26__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_28__pin_a2f_o_1_, chanx_left_in[93]}),
		.sram(mux_tree_tapbuf_L4SB_size13_8_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size13_8_sram_inv[0:3]),
		.out(chany_bottom_out[92]));

	mux_tree_tapbuf_L4SB_size13 mux_bottom_track_189 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_25__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_27__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_29__pin_a2f_o_1_, chanx_left_in[95]}),
		.sram(mux_tree_tapbuf_L4SB_size13_9_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size13_9_sram_inv[0:3]),
		.out(chany_bottom_out[94]));

	mux_tree_tapbuf_L4SB_size13 mux_left_track_39 (
		.in({chany_bottom_in[18], left_bottom_grid_top_width_0_height_0_subtile_30__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_32__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_36__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_37__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_40__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_44__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_44__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_48__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_51__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_52__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_56__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_58__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size13_10_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size13_10_sram_inv[0:3]),
		.out(chanx_left_out[19]));

	mux_tree_tapbuf_L4SB_size13 mux_left_track_43 (
		.in({chany_bottom_in[20], left_bottom_grid_top_width_0_height_0_subtile_31__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_33__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_37__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_38__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_41__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_45__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_45__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_49__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_52__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_53__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_57__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_59__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size13_11_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size13_11_sram_inv[0:3]),
		.out(chanx_left_out[21]));

	mux_tree_tapbuf_L4SB_size13 mux_left_track_137 (
		.in({chany_bottom_in[67], left_bottom_grid_top_width_0_height_0_subtile_30__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_30__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_34__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_37__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_38__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_42__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_44__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_46__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_50__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_51__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_54__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_58__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size13_12_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size13_12_sram_inv[0:3]),
		.out(chanx_left_out[68]));

	mux_tree_tapbuf_L4SB_size13 mux_left_track_141 (
		.in({chany_bottom_in[69], left_bottom_grid_top_width_0_height_0_subtile_31__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_31__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_35__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_38__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_39__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_43__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_45__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_47__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_51__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_52__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_55__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_59__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size13_13_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size13_13_sram_inv[0:3]),
		.out(chanx_left_out[70]));

	mux_tree_tapbuf_L4SB_size13 mux_left_track_153 (
		.in({chany_bottom_in[75], left_bottom_grid_top_width_0_height_0_subtile_30__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_34__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_34__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_38__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_41__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_42__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_46__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_48__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_50__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_54__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_55__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_58__pin_a2f_o_1_}),
		.sram(mux_tree_tapbuf_L4SB_size13_14_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size13_14_sram_inv[0:3]),
		.out(chanx_left_out[76]));

	mux_tree_tapbuf_L4SB_size13 mux_left_track_157 (
		.in({chany_bottom_in[77], left_bottom_grid_top_width_0_height_0_subtile_31__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_35__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_35__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_39__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_42__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_43__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_47__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_49__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_51__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_55__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_56__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_59__pin_a2f_o_1_}),
		.sram(mux_tree_tapbuf_L4SB_size13_15_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size13_15_sram_inv[0:3]),
		.out(chanx_left_out[78]));

	mux_tree_tapbuf_L4SB_size13 mux_left_track_165 (
		.in({chany_bottom_in[81], left_bottom_grid_top_width_0_height_0_subtile_30__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_33__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_37__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_37__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_41__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_44__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_45__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_49__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_51__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_53__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_57__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_58__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size13_16_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size13_16_sram_inv[0:3]),
		.out(chanx_left_out[82]));

	mux_tree_tapbuf_L4SB_size13 mux_left_track_173 (
		.in({chany_bottom_in[85], left_bottom_grid_top_width_0_height_0_subtile_31__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_32__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_35__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_39__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_39__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_43__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_46__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_47__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_51__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_53__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_55__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_59__pin_a2f_o_1_}),
		.sram(mux_tree_tapbuf_L4SB_size13_17_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size13_17_sram_inv[0:3]),
		.out(chanx_left_out[86]));

	mux_tree_tapbuf_L4SB_size13 mux_left_track_185 (
		.in({chany_bottom_in[91], left_bottom_grid_top_width_0_height_0_subtile_30__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_34__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_35__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_38__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_42__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_42__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_46__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_49__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_50__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_54__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_56__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_58__pin_a2f_o_1_}),
		.sram(mux_tree_tapbuf_L4SB_size13_18_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size13_18_sram_inv[0:3]),
		.out(chanx_left_out[92]));

	mux_tree_tapbuf_L4SB_size13 mux_left_track_189 (
		.in({chany_bottom_in[93], left_bottom_grid_top_width_0_height_0_subtile_31__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_35__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_36__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_39__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_43__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_43__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_47__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_50__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_51__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_55__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_57__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_59__pin_a2f_o_1_}),
		.sram(mux_tree_tapbuf_L4SB_size13_19_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size13_19_sram_inv[0:3]),
		.out(chanx_left_out[94]));

	mux_tree_tapbuf_L4SB_size13_mem mem_bottom_track_39 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size13_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size13_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size13_0_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size13_mem mem_bottom_track_43 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size6_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size13_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size13_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size13_1_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size13_mem mem_bottom_track_137 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size6_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size13_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size13_2_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size13_2_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size13_mem mem_bottom_track_141 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size6_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size13_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size13_3_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size13_3_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size13_mem mem_bottom_track_153 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size6_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size13_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size13_4_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size13_4_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size13_mem mem_bottom_track_157 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size6_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size13_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size13_5_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size13_5_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size13_mem mem_bottom_track_165 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size5_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size13_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size13_6_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size13_6_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size13_mem mem_bottom_track_173 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size5_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size13_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size13_7_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size13_7_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size13_mem mem_bottom_track_185 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size6_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size13_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size13_8_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size13_8_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size13_mem mem_bottom_track_189 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size5_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size13_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size13_9_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size13_9_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size13_mem mem_left_track_39 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_31_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size13_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size13_10_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size13_10_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size13_mem mem_left_track_43 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size6_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size13_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size13_11_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size13_11_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size13_mem mem_left_track_137 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size6_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size13_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size13_12_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size13_12_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size13_mem mem_left_track_141 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size6_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size13_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size13_13_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size13_13_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size13_mem mem_left_track_153 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size6_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size13_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size13_14_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size13_14_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size13_mem mem_left_track_157 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size6_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size13_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size13_15_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size13_15_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size13_mem mem_left_track_165 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size5_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size13_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size13_16_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size13_16_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size13_mem mem_left_track_173 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size5_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size13_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size13_17_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size13_17_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size13_mem mem_left_track_185 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size6_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size13_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size13_18_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size13_18_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size13_mem mem_left_track_189 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size5_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size13_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size13_19_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size13_19_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size6 mux_bottom_track_41 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_25__pin_a2f_o_0_, chanx_left_in[21]}),
		.sram(mux_tree_tapbuf_L4SB_size6_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size6_0_sram_inv[0:2]),
		.out(chany_bottom_out[20]));

	mux_tree_tapbuf_L4SB_size6 mux_bottom_track_45 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_26__pin_a2f_o_0_, chanx_left_in[23]}),
		.sram(mux_tree_tapbuf_L4SB_size6_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size6_1_sram_inv[0:2]),
		.out(chany_bottom_out[22]));

	mux_tree_tapbuf_L4SB_size6 mux_bottom_track_49 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_27__pin_a2f_o_0_, chanx_left_in[25]}),
		.sram(mux_tree_tapbuf_L4SB_size6_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size6_2_sram_inv[0:2]),
		.out(chany_bottom_out[24]));

	mux_tree_tapbuf_L4SB_size6 mux_bottom_track_135 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_24__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_26__pin_a2f_o_1_, chanx_left_in[68]}),
		.sram(mux_tree_tapbuf_L4SB_size6_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size6_3_sram_inv[0:2]),
		.out(chany_bottom_out[67]));

	mux_tree_tapbuf_L4SB_size6 mux_bottom_track_139 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_25__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_27__pin_a2f_o_1_, chanx_left_in[70]}),
		.sram(mux_tree_tapbuf_L4SB_size6_4_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size6_4_sram_inv[0:2]),
		.out(chany_bottom_out[69]));

	mux_tree_tapbuf_L4SB_size6 mux_bottom_track_143 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_26__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_28__pin_a2f_o_1_, chanx_left_in[72]}),
		.sram(mux_tree_tapbuf_L4SB_size6_5_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size6_5_sram_inv[0:2]),
		.out(chany_bottom_out[71]));

	mux_tree_tapbuf_L4SB_size6 mux_bottom_track_147 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_27__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_29__pin_a2f_o_1_, chanx_left_in[74]}),
		.sram(mux_tree_tapbuf_L4SB_size6_6_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size6_6_sram_inv[0:2]),
		.out(chany_bottom_out[73]));

	mux_tree_tapbuf_L4SB_size6 mux_bottom_track_151 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_28__pin_a2f_o_0_, chanx_left_in[76]}),
		.sram(mux_tree_tapbuf_L4SB_size6_7_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size6_7_sram_inv[0:2]),
		.out(chany_bottom_out[75]));

	mux_tree_tapbuf_L4SB_size6 mux_bottom_track_155 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_29__pin_a2f_o_0_, chanx_left_in[78]}),
		.sram(mux_tree_tapbuf_L4SB_size6_8_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size6_8_sram_inv[0:2]),
		.out(chany_bottom_out[77]));

	mux_tree_tapbuf_L4SB_size6 mux_bottom_track_179 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_28__pin_a2f_o_0_, chanx_left_in[90]}),
		.sram(mux_tree_tapbuf_L4SB_size6_9_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size6_9_sram_inv[0:2]),
		.out(chany_bottom_out[89]));

	mux_tree_tapbuf_L4SB_size6 mux_bottom_track_183 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_29__pin_a2f_o_0_, chanx_left_in[92]}),
		.sram(mux_tree_tapbuf_L4SB_size6_10_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size6_10_sram_inv[0:2]),
		.out(chany_bottom_out[91]));

	mux_tree_tapbuf_L4SB_size6 mux_left_track_41 (
		.in({chany_bottom_in[19], left_bottom_grid_top_width_0_height_0_subtile_30__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_34__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_41__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_48__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_55__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size6_11_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size6_11_sram_inv[0:2]),
		.out(chanx_left_out[20]));

	mux_tree_tapbuf_L4SB_size6 mux_left_track_45 (
		.in({chany_bottom_in[21], left_bottom_grid_top_width_0_height_0_subtile_31__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_35__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_42__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_49__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_56__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size6_12_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size6_12_sram_inv[0:2]),
		.out(chanx_left_out[22]));

	mux_tree_tapbuf_L4SB_size6 mux_left_track_49 (
		.in({chany_bottom_in[23], left_bottom_grid_top_width_0_height_0_subtile_32__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_36__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_43__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_50__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_57__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size6_13_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size6_13_sram_inv[0:2]),
		.out(chanx_left_out[24]));

	mux_tree_tapbuf_L4SB_size6 mux_left_track_135 (
		.in({chany_bottom_in[66], left_bottom_grid_top_width_0_height_0_subtile_33__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_40__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_47__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_54__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_56__pin_a2f_o_1_}),
		.sram(mux_tree_tapbuf_L4SB_size6_14_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size6_14_sram_inv[0:2]),
		.out(chanx_left_out[67]));

	mux_tree_tapbuf_L4SB_size6 mux_left_track_139 (
		.in({chany_bottom_in[68], left_bottom_grid_top_width_0_height_0_subtile_34__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_41__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_48__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_55__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_57__pin_a2f_o_1_}),
		.sram(mux_tree_tapbuf_L4SB_size6_15_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size6_15_sram_inv[0:2]),
		.out(chanx_left_out[69]));

	mux_tree_tapbuf_L4SB_size6 mux_left_track_143 (
		.in({chany_bottom_in[70], left_bottom_grid_top_width_0_height_0_subtile_35__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_42__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_49__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_56__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_58__pin_a2f_o_1_}),
		.sram(mux_tree_tapbuf_L4SB_size6_16_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size6_16_sram_inv[0:2]),
		.out(chanx_left_out[71]));

	mux_tree_tapbuf_L4SB_size6 mux_left_track_147 (
		.in({chany_bottom_in[72], left_bottom_grid_top_width_0_height_0_subtile_36__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_43__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_50__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_57__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_59__pin_a2f_o_1_}),
		.sram(mux_tree_tapbuf_L4SB_size6_17_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size6_17_sram_inv[0:2]),
		.out(chanx_left_out[73]));

	mux_tree_tapbuf_L4SB_size6 mux_left_track_151 (
		.in({chany_bottom_in[74], left_bottom_grid_top_width_0_height_0_subtile_30__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_37__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_44__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_51__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_58__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size6_18_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size6_18_sram_inv[0:2]),
		.out(chanx_left_out[75]));

	mux_tree_tapbuf_L4SB_size6 mux_left_track_155 (
		.in({chany_bottom_in[76], left_bottom_grid_top_width_0_height_0_subtile_31__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_38__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_45__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_52__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_59__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size6_19_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size6_19_sram_inv[0:2]),
		.out(chanx_left_out[77]));

	mux_tree_tapbuf_L4SB_size6 mux_left_track_179 (
		.in({chany_bottom_in[88], left_bottom_grid_top_width_0_height_0_subtile_30__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_37__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_44__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_51__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_58__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size6_20_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size6_20_sram_inv[0:2]),
		.out(chanx_left_out[89]));

	mux_tree_tapbuf_L4SB_size6 mux_left_track_183 (
		.in({chany_bottom_in[90], left_bottom_grid_top_width_0_height_0_subtile_31__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_38__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_45__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_52__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_59__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size6_21_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size6_21_sram_inv[0:2]),
		.out(chanx_left_out[91]));

	mux_tree_tapbuf_L4SB_size6_mem mem_bottom_track_41 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size13_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size6_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size6_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size6_0_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size6_mem mem_bottom_track_45 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size13_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size6_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size6_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size6_1_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size6_mem mem_bottom_track_49 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size12_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size6_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size6_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size6_2_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size6_mem mem_bottom_track_135 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size11_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size6_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size6_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size6_3_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size6_mem mem_bottom_track_139 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size13_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size6_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size6_4_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size6_4_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size6_mem mem_bottom_track_143 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size13_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size6_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size6_5_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size6_5_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size6_mem mem_bottom_track_147 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size12_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size6_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size6_6_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size6_6_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size6_mem mem_bottom_track_151 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size12_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size6_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size6_7_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size6_7_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size6_mem mem_bottom_track_155 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size13_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size6_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size6_8_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size6_8_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size6_mem mem_bottom_track_179 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size12_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size6_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size6_9_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size6_9_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size6_mem mem_bottom_track_183 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size12_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size6_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size6_10_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size6_10_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size6_mem mem_left_track_41 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size13_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size6_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size6_11_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size6_11_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size6_mem mem_left_track_45 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size13_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size6_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size6_12_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size6_12_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size6_mem mem_left_track_49 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size12_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size6_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size6_13_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size6_13_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size6_mem mem_left_track_135 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size11_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size6_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size6_14_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size6_14_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size6_mem mem_left_track_139 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size13_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size6_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size6_15_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size6_15_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size6_mem mem_left_track_143 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size13_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size6_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size6_16_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size6_16_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size6_mem mem_left_track_147 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size12_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size6_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size6_17_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size6_17_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size6_mem mem_left_track_151 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size12_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size6_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size6_18_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size6_18_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size6_mem mem_left_track_155 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size13_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size6_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size6_19_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size6_19_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size6_mem mem_left_track_179 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size12_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size6_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size6_20_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size6_20_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size6_mem mem_left_track_183 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size12_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size6_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size6_21_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size6_21_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size12 mux_bottom_track_47 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_24__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_28__pin_a2f_o_1_, chanx_left_in[24]}),
		.sram(mux_tree_tapbuf_L4SB_size12_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size12_0_sram_inv[0:3]),
		.out(chany_bottom_out[23]));

	mux_tree_tapbuf_L4SB_size12 mux_bottom_track_51 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_24__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_25__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_29__pin_a2f_o_1_, chanx_left_in[26]}),
		.sram(mux_tree_tapbuf_L4SB_size12_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size12_1_sram_inv[0:3]),
		.out(chany_bottom_out[25]));

	mux_tree_tapbuf_L4SB_size12 mux_bottom_track_67 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_25__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_28__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_29__pin_a2f_o_1_, chanx_left_in[34]}),
		.sram(mux_tree_tapbuf_L4SB_size12_2_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size12_2_sram_inv[0:3]),
		.out(chany_bottom_out[33]));

	mux_tree_tapbuf_L4SB_size12 mux_bottom_track_145 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_26__pin_a2f_o_1_, chanx_left_in[73]}),
		.sram(mux_tree_tapbuf_L4SB_size12_3_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size12_3_sram_inv[0:3]),
		.out(chany_bottom_out[72]));

	mux_tree_tapbuf_L4SB_size12 mux_bottom_track_149 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_24__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_27__pin_a2f_o_1_, chanx_left_in[75]}),
		.sram(mux_tree_tapbuf_L4SB_size12_4_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size12_4_sram_inv[0:3]),
		.out(chany_bottom_out[74]));

	mux_tree_tapbuf_L4SB_size12 mux_bottom_track_161 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_26__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_27__pin_a2f_o_0_, chanx_left_in[81]}),
		.sram(mux_tree_tapbuf_L4SB_size12_5_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size12_5_sram_inv[0:3]),
		.out(chany_bottom_out[80]));

	mux_tree_tapbuf_L4SB_size12 mux_bottom_track_177 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_24__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_26__pin_a2f_o_1_, chanx_left_in[89]}),
		.sram(mux_tree_tapbuf_L4SB_size12_6_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size12_6_sram_inv[0:3]),
		.out(chany_bottom_out[88]));

	mux_tree_tapbuf_L4SB_size12 mux_bottom_track_181 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_25__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_27__pin_a2f_o_1_, chanx_left_in[91]}),
		.sram(mux_tree_tapbuf_L4SB_size12_7_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size12_7_sram_inv[0:3]),
		.out(chany_bottom_out[90]));

	mux_tree_tapbuf_L4SB_size12 mux_left_track_47 (
		.in({chany_bottom_in[22], left_bottom_grid_top_width_0_height_0_subtile_32__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_34__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_38__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_39__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_42__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_46__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_46__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_50__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_53__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_54__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_58__pin_a2f_o_1_}),
		.sram(mux_tree_tapbuf_L4SB_size12_8_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size12_8_sram_inv[0:3]),
		.out(chanx_left_out[23]));

	mux_tree_tapbuf_L4SB_size12 mux_left_track_51 (
		.in({chany_bottom_in[24], left_bottom_grid_top_width_0_height_0_subtile_33__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_35__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_39__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_40__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_43__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_47__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_47__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_51__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_54__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_55__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_59__pin_a2f_o_1_}),
		.sram(mux_tree_tapbuf_L4SB_size12_9_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size12_9_sram_inv[0:3]),
		.out(chanx_left_out[25]));

	mux_tree_tapbuf_L4SB_size12 mux_left_track_67 (
		.in({chany_bottom_in[32], left_bottom_grid_top_width_0_height_0_subtile_30__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_37__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_39__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_43__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_44__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_47__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_51__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_51__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_55__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_58__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_59__pin_a2f_o_1_}),
		.sram(mux_tree_tapbuf_L4SB_size12_10_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size12_10_sram_inv[0:3]),
		.out(chanx_left_out[33]));

	mux_tree_tapbuf_L4SB_size12 mux_left_track_145 (
		.in({chany_bottom_in[71], left_bottom_grid_top_width_0_height_0_subtile_32__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_32__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_36__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_39__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_40__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_44__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_46__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_48__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_52__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_53__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_56__pin_a2f_o_1_}),
		.sram(mux_tree_tapbuf_L4SB_size12_11_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size12_11_sram_inv[0:3]),
		.out(chanx_left_out[72]));

	mux_tree_tapbuf_L4SB_size12 mux_left_track_149 (
		.in({chany_bottom_in[73], left_bottom_grid_top_width_0_height_0_subtile_33__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_33__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_37__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_40__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_41__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_45__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_47__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_49__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_53__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_54__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_57__pin_a2f_o_1_}),
		.sram(mux_tree_tapbuf_L4SB_size12_12_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size12_12_sram_inv[0:3]),
		.out(chanx_left_out[74]));

	mux_tree_tapbuf_L4SB_size12 mux_left_track_161 (
		.in({chany_bottom_in[79], left_bottom_grid_top_width_0_height_0_subtile_32__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_36__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_36__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_40__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_43__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_44__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_48__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_50__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_52__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_56__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_57__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size12_13_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size12_13_sram_inv[0:3]),
		.out(chanx_left_out[80]));

	mux_tree_tapbuf_L4SB_size12 mux_left_track_177 (
		.in({chany_bottom_in[87], left_bottom_grid_top_width_0_height_0_subtile_32__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_33__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_36__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_40__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_40__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_44__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_47__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_48__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_52__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_54__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_56__pin_a2f_o_1_}),
		.sram(mux_tree_tapbuf_L4SB_size12_14_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size12_14_sram_inv[0:3]),
		.out(chanx_left_out[88]));

	mux_tree_tapbuf_L4SB_size12 mux_left_track_181 (
		.in({chany_bottom_in[89], left_bottom_grid_top_width_0_height_0_subtile_33__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_34__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_37__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_41__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_41__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_45__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_48__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_49__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_53__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_55__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_57__pin_a2f_o_1_}),
		.sram(mux_tree_tapbuf_L4SB_size12_15_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size12_15_sram_inv[0:3]),
		.out(chanx_left_out[90]));

	mux_tree_tapbuf_L4SB_size12_mem mem_bottom_track_47 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size6_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size12_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size12_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size12_0_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size12_mem mem_bottom_track_51 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size6_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size12_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size12_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size12_1_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size12_mem mem_bottom_track_67 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size7_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size12_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size12_2_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size12_2_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size12_mem mem_bottom_track_145 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size6_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size12_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size12_3_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size12_3_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size12_mem mem_bottom_track_149 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size6_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size12_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size12_4_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size12_4_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size12_mem mem_bottom_track_161 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size5_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size12_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size12_5_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size12_5_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size12_mem mem_bottom_track_177 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size5_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size12_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size12_6_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size12_6_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size12_mem mem_bottom_track_181 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size6_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size12_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size12_7_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size12_7_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size12_mem mem_left_track_47 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size6_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size12_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size12_8_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size12_8_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size12_mem mem_left_track_51 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size6_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size12_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size12_9_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size12_9_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size12_mem mem_left_track_67 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size7_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size12_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size12_10_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size12_10_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size12_mem mem_left_track_145 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size6_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size12_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size12_11_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size12_11_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size12_mem mem_left_track_149 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size6_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size12_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size12_12_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size12_12_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size12_mem mem_left_track_161 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size5_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size12_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size12_13_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size12_13_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size12_mem mem_left_track_177 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size5_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size12_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size12_14_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size12_14_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size12_mem mem_left_track_181 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size6_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size12_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size12_15_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size12_15_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size7 mux_bottom_track_53 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_28__pin_a2f_o_0_, chanx_left_in[27]}),
		.sram(mux_tree_tapbuf_L4SB_size7_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_0_sram_inv[0:2]),
		.out(chany_bottom_out[26]));

	mux_tree_tapbuf_L4SB_size7 mux_bottom_track_61 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_, chanx_left_in[31]}),
		.sram(mux_tree_tapbuf_L4SB_size7_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_1_sram_inv[0:2]),
		.out(chany_bottom_out[30]));

	mux_tree_tapbuf_L4SB_size7 mux_bottom_track_65 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_24__pin_a2f_o_0_, chanx_left_in[33]}),
		.sram(mux_tree_tapbuf_L4SB_size7_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_2_sram_inv[0:2]),
		.out(chany_bottom_out[32]));

	mux_tree_tapbuf_L4SB_size7 mux_bottom_track_69 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_25__pin_a2f_o_0_, chanx_left_in[35]}),
		.sram(mux_tree_tapbuf_L4SB_size7_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_3_sram_inv[0:2]),
		.out(chany_bottom_out[34]));

	mux_tree_tapbuf_L4SB_size7 mux_bottom_track_119 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_26__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_27__pin_a2f_o_0_, chanx_left_in[60]}),
		.sram(mux_tree_tapbuf_L4SB_size7_4_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_4_sram_inv[0:2]),
		.out(chany_bottom_out[59]));

	mux_tree_tapbuf_L4SB_size7 mux_bottom_track_131 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_25__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_29__pin_a2f_o_1_, chanx_left_in[66]}),
		.sram(mux_tree_tapbuf_L4SB_size7_5_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_5_sram_inv[0:2]),
		.out(chany_bottom_out[65]));

	mux_tree_tapbuf_L4SB_size7 mux_left_track_53 (
		.in({chany_bottom_in[25], left_bottom_grid_top_width_0_height_0_subtile_30__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_33__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_37__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_44__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_51__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_58__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size7_6_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_6_sram_inv[0:2]),
		.out(chanx_left_out[26]));

	mux_tree_tapbuf_L4SB_size7 mux_left_track_61 (
		.in({chany_bottom_in[29], left_bottom_grid_top_width_0_height_0_subtile_31__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_32__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_35__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_39__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_46__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_53__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size7_7_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_7_sram_inv[0:2]),
		.out(chanx_left_out[30]));

	mux_tree_tapbuf_L4SB_size7 mux_left_track_65 (
		.in({chany_bottom_in[31], left_bottom_grid_top_width_0_height_0_subtile_32__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_33__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_36__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_40__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_47__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_54__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size7_8_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_8_sram_inv[0:2]),
		.out(chanx_left_out[32]));

	mux_tree_tapbuf_L4SB_size7 mux_left_track_69 (
		.in({chany_bottom_in[33], left_bottom_grid_top_width_0_height_0_subtile_33__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_34__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_37__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_41__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_48__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_55__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size7_9_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_9_sram_inv[0:2]),
		.out(chanx_left_out[34]));

	mux_tree_tapbuf_L4SB_size7 mux_left_track_119 (
		.in({chany_bottom_in[58], left_bottom_grid_top_width_0_height_0_subtile_36__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_43__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_50__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_52__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_56__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_57__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size7_10_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_10_sram_inv[0:2]),
		.out(chanx_left_out[59]));

	mux_tree_tapbuf_L4SB_size7 mux_left_track_131 (
		.in({chany_bottom_in[64], left_bottom_grid_top_width_0_height_0_subtile_32__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_39__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_46__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_53__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_55__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_59__pin_a2f_o_1_}),
		.sram(mux_tree_tapbuf_L4SB_size7_11_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_11_sram_inv[0:2]),
		.out(chanx_left_out[65]));

	mux_tree_tapbuf_L4SB_size7_mem mem_bottom_track_53 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size12_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size7_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size7_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_0_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7_mem mem_bottom_track_61 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size11_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size7_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size7_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_1_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7_mem mem_bottom_track_65 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size11_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size7_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size7_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_2_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7_mem mem_bottom_track_69 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size12_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size7_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size7_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_3_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7_mem mem_bottom_track_119 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size10_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size7_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size7_4_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_4_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7_mem mem_bottom_track_131 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size11_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size7_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size7_5_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_5_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7_mem mem_left_track_53 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size12_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size7_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size7_6_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_6_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7_mem mem_left_track_61 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size11_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size7_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size7_7_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_7_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7_mem mem_left_track_65 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size11_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size7_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size7_8_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_8_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7_mem mem_left_track_69 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size12_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size7_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size7_9_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_9_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7_mem mem_left_track_119 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size10_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size7_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size7_10_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_10_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7_mem mem_left_track_131 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size11_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size7_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size7_11_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_11_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size11 mux_bottom_track_55 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_25__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_26__pin_a2f_o_1_, chanx_left_in[28]}),
		.sram(mux_tree_tapbuf_L4SB_size11_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size11_0_sram_inv[0:3]),
		.out(chany_bottom_out[27]));

	mux_tree_tapbuf_L4SB_size11 mux_bottom_track_59 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_26__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_27__pin_a2f_o_1_, chanx_left_in[30]}),
		.sram(mux_tree_tapbuf_L4SB_size11_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size11_1_sram_inv[0:3]),
		.out(chany_bottom_out[29]));

	mux_tree_tapbuf_L4SB_size11 mux_bottom_track_63 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_24__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_27__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_28__pin_a2f_o_1_, chanx_left_in[32]}),
		.sram(mux_tree_tapbuf_L4SB_size11_2_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size11_2_sram_inv[0:3]),
		.out(chany_bottom_out[31]));

	mux_tree_tapbuf_L4SB_size11 mux_bottom_track_71 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_26__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_29__pin_a2f_o_0_, chanx_left_in[36]}),
		.sram(mux_tree_tapbuf_L4SB_size11_3_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size11_3_sram_inv[0:3]),
		.out(chany_bottom_out[35]));

	mux_tree_tapbuf_L4SB_size11 mux_bottom_track_109 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_28__pin_a2f_o_0_, chanx_left_in[55]}),
		.sram(mux_tree_tapbuf_L4SB_size11_4_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size11_4_sram_inv[0:3]),
		.out(chany_bottom_out[54]));

	mux_tree_tapbuf_L4SB_size11 mux_bottom_track_113 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_29__pin_a2f_o_0_, chanx_left_in[57]}),
		.sram(mux_tree_tapbuf_L4SB_size11_5_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size11_5_sram_inv[0:3]),
		.out(chany_bottom_out[56]));

	mux_tree_tapbuf_L4SB_size11 mux_bottom_track_121 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_24__pin_a2f_o_0_, chanx_left_in[61]}),
		.sram(mux_tree_tapbuf_L4SB_size11_6_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size11_6_sram_inv[0:3]),
		.out(chany_bottom_out[60]));

	mux_tree_tapbuf_L4SB_size11 mux_bottom_track_125 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_25__pin_a2f_o_0_, chanx_left_in[63]}),
		.sram(mux_tree_tapbuf_L4SB_size11_7_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size11_7_sram_inv[0:3]),
		.out(chany_bottom_out[62]));

	mux_tree_tapbuf_L4SB_size11 mux_bottom_track_129 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_26__pin_a2f_o_0_, chanx_left_in[65]}),
		.sram(mux_tree_tapbuf_L4SB_size11_8_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size11_8_sram_inv[0:3]),
		.out(chany_bottom_out[64]));

	mux_tree_tapbuf_L4SB_size11 mux_bottom_track_133 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_27__pin_a2f_o_0_, chanx_left_in[67]}),
		.sram(mux_tree_tapbuf_L4SB_size11_9_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size11_9_sram_inv[0:3]),
		.out(chany_bottom_out[66]));

	mux_tree_tapbuf_L4SB_size11 mux_left_track_55 (
		.in({chany_bottom_in[26], left_bottom_grid_top_width_0_height_0_subtile_34__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_36__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_40__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_41__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_44__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_48__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_48__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_52__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_55__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_56__pin_a2f_o_1_}),
		.sram(mux_tree_tapbuf_L4SB_size11_10_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size11_10_sram_inv[0:3]),
		.out(chanx_left_out[27]));

	mux_tree_tapbuf_L4SB_size11 mux_left_track_59 (
		.in({chany_bottom_in[28], left_bottom_grid_top_width_0_height_0_subtile_35__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_37__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_41__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_42__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_45__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_49__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_49__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_53__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_56__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_57__pin_a2f_o_1_}),
		.sram(mux_tree_tapbuf_L4SB_size11_11_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size11_11_sram_inv[0:3]),
		.out(chanx_left_out[29]));

	mux_tree_tapbuf_L4SB_size11 mux_left_track_63 (
		.in({chany_bottom_in[30], left_bottom_grid_top_width_0_height_0_subtile_36__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_38__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_42__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_43__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_46__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_50__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_50__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_54__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_57__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_58__pin_a2f_o_1_}),
		.sram(mux_tree_tapbuf_L4SB_size11_12_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size11_12_sram_inv[0:3]),
		.out(chanx_left_out[31]));

	mux_tree_tapbuf_L4SB_size11 mux_left_track_71 (
		.in({chany_bottom_in[34], left_bottom_grid_top_width_0_height_0_subtile_31__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_38__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_40__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_44__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_45__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_48__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_52__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_52__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_56__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_59__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size11_13_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size11_13_sram_inv[0:3]),
		.out(chanx_left_out[35]));

	mux_tree_tapbuf_L4SB_size11 mux_left_track_109 (
		.in({chany_bottom_in[53], left_bottom_grid_top_width_0_height_0_subtile_30__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_31__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_35__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_37__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_39__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_43__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_44__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_47__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_51__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_58__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size11_14_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size11_14_sram_inv[0:3]),
		.out(chanx_left_out[54]));

	mux_tree_tapbuf_L4SB_size11 mux_left_track_113 (
		.in({chany_bottom_in[55], left_bottom_grid_top_width_0_height_0_subtile_31__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_32__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_36__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_38__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_40__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_44__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_45__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_48__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_52__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_59__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size11_15_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size11_15_sram_inv[0:3]),
		.out(chanx_left_out[56]));

	mux_tree_tapbuf_L4SB_size11 mux_left_track_121 (
		.in({chany_bottom_in[59], left_bottom_grid_top_width_0_height_0_subtile_30__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_33__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_34__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_38__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_40__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_42__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_46__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_47__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_50__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_54__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size11_16_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size11_16_sram_inv[0:3]),
		.out(chanx_left_out[60]));

	mux_tree_tapbuf_L4SB_size11 mux_left_track_125 (
		.in({chany_bottom_in[61], left_bottom_grid_top_width_0_height_0_subtile_31__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_34__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_35__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_39__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_41__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_43__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_47__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_48__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_51__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_55__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size11_17_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size11_17_sram_inv[0:3]),
		.out(chanx_left_out[62]));

	mux_tree_tapbuf_L4SB_size11 mux_left_track_129 (
		.in({chany_bottom_in[63], left_bottom_grid_top_width_0_height_0_subtile_32__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_35__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_36__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_40__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_42__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_44__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_48__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_49__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_52__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_56__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size11_18_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size11_18_sram_inv[0:3]),
		.out(chanx_left_out[64]));

	mux_tree_tapbuf_L4SB_size11 mux_left_track_133 (
		.in({chany_bottom_in[65], left_bottom_grid_top_width_0_height_0_subtile_33__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_36__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_37__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_41__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_43__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_45__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_49__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_50__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_53__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_57__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size11_19_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size11_19_sram_inv[0:3]),
		.out(chanx_left_out[66]));

	mux_tree_tapbuf_L4SB_size11_mem mem_bottom_track_55 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size7_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size11_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size11_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size11_0_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size11_mem mem_bottom_track_59 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size11_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size11_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size11_1_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size11_mem mem_bottom_track_63 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size7_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size11_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size11_2_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size11_2_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size11_mem mem_bottom_track_71 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size7_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size11_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size11_3_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size11_3_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size11_mem mem_bottom_track_109 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size11_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size11_4_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size11_4_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size11_mem mem_bottom_track_113 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size11_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size11_5_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size11_5_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size11_mem mem_bottom_track_121 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size7_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size11_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size11_6_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size11_6_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size11_mem mem_bottom_track_125 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size11_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size11_7_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size11_7_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size11_mem mem_bottom_track_129 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size11_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size11_8_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size11_8_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size11_mem mem_bottom_track_133 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size7_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size11_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size11_9_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size11_9_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size11_mem mem_left_track_55 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size7_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size11_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size11_10_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size11_10_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size11_mem mem_left_track_59 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size11_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size11_11_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size11_11_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size11_mem mem_left_track_63 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size7_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size11_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size11_12_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size11_12_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size11_mem mem_left_track_71 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size7_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size11_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size11_13_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size11_13_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size11_mem mem_left_track_109 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size11_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size11_14_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size11_14_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size11_mem mem_left_track_113 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size11_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size11_15_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size11_15_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size11_mem mem_left_track_121 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size7_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size11_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size11_16_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size11_16_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size11_mem mem_left_track_125 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size11_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size11_17_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size11_17_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size11_mem mem_left_track_129 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size11_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size11_18_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size11_18_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size11_mem mem_left_track_133 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size7_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size11_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size11_19_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size11_19_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_57 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_29__pin_a2f_o_0_, chanx_left_in[29]}),
		.sram(mux_tree_tapbuf_L4SB_size8_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_0_sram_inv[0:2]),
		.out(chany_bottom_out[28]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_73 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_26__pin_a2f_o_0_, chanx_left_in[37]}),
		.sram(mux_tree_tapbuf_L4SB_size8_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_1_sram_inv[0:2]),
		.out(chany_bottom_out[36]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_77 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_27__pin_a2f_o_0_, chanx_left_in[39]}),
		.sram(mux_tree_tapbuf_L4SB_size8_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_2_sram_inv[0:2]),
		.out(chany_bottom_out[38]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_103 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_26__pin_a2f_o_1_, chanx_left_in[52]}),
		.sram(mux_tree_tapbuf_L4SB_size8_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_3_sram_inv[0:2]),
		.out(chany_bottom_out[51]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_107 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_24__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_27__pin_a2f_o_1_, chanx_left_in[54]}),
		.sram(mux_tree_tapbuf_L4SB_size8_4_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_4_sram_inv[0:2]),
		.out(chany_bottom_out[53]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_111 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_24__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_25__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_28__pin_a2f_o_1_, chanx_left_in[56]}),
		.sram(mux_tree_tapbuf_L4SB_size8_5_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_5_sram_inv[0:2]),
		.out(chany_bottom_out[55]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_115 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_25__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_26__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_29__pin_a2f_o_1_, chanx_left_in[58]}),
		.sram(mux_tree_tapbuf_L4SB_size8_6_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_6_sram_inv[0:2]),
		.out(chany_bottom_out[57]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_123 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_27__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_28__pin_a2f_o_0_, chanx_left_in[62]}),
		.sram(mux_tree_tapbuf_L4SB_size8_7_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_7_sram_inv[0:2]),
		.out(chany_bottom_out[61]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_127 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_24__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_28__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_29__pin_a2f_o_0_, chanx_left_in[64]}),
		.sram(mux_tree_tapbuf_L4SB_size8_8_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_8_sram_inv[0:2]),
		.out(chany_bottom_out[63]));

	mux_tree_tapbuf_L4SB_size8 mux_left_track_57 (
		.in({chany_bottom_in[27], left_bottom_grid_top_width_0_height_0_subtile_30__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_31__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_34__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_38__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_45__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_52__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_59__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_9_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_9_sram_inv[0:2]),
		.out(chanx_left_out[28]));

	mux_tree_tapbuf_L4SB_size8 mux_left_track_73 (
		.in({chany_bottom_in[35], left_bottom_grid_top_width_0_height_0_subtile_30__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_34__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_35__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_38__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_42__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_49__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_56__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_10_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_10_sram_inv[0:2]),
		.out(chanx_left_out[36]));

	mux_tree_tapbuf_L4SB_size8 mux_left_track_77 (
		.in({chany_bottom_in[37], left_bottom_grid_top_width_0_height_0_subtile_31__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_35__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_36__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_39__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_43__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_50__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_57__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_11_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_11_sram_inv[0:2]),
		.out(chanx_left_out[38]));

	mux_tree_tapbuf_L4SB_size8 mux_left_track_103 (
		.in({chany_bottom_in[50], left_bottom_grid_top_width_0_height_0_subtile_32__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_39__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_46__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_48__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_52__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_53__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_56__pin_a2f_o_1_}),
		.sram(mux_tree_tapbuf_L4SB_size8_12_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_12_sram_inv[0:2]),
		.out(chanx_left_out[51]));

	mux_tree_tapbuf_L4SB_size8 mux_left_track_107 (
		.in({chany_bottom_in[52], left_bottom_grid_top_width_0_height_0_subtile_33__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_40__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_47__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_49__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_53__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_54__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_57__pin_a2f_o_1_}),
		.sram(mux_tree_tapbuf_L4SB_size8_13_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_13_sram_inv[0:2]),
		.out(chanx_left_out[53]));

	mux_tree_tapbuf_L4SB_size8 mux_left_track_111 (
		.in({chany_bottom_in[54], left_bottom_grid_top_width_0_height_0_subtile_34__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_41__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_48__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_50__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_54__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_55__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_58__pin_a2f_o_1_}),
		.sram(mux_tree_tapbuf_L4SB_size8_14_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_14_sram_inv[0:2]),
		.out(chanx_left_out[55]));

	mux_tree_tapbuf_L4SB_size8 mux_left_track_115 (
		.in({chany_bottom_in[56], left_bottom_grid_top_width_0_height_0_subtile_35__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_42__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_49__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_51__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_55__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_56__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_59__pin_a2f_o_1_}),
		.sram(mux_tree_tapbuf_L4SB_size8_15_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_15_sram_inv[0:2]),
		.out(chanx_left_out[57]));

	mux_tree_tapbuf_L4SB_size8 mux_left_track_123 (
		.in({chany_bottom_in[60], left_bottom_grid_top_width_0_height_0_subtile_30__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_37__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_44__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_51__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_53__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_57__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_58__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_16_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_16_sram_inv[0:2]),
		.out(chanx_left_out[61]));

	mux_tree_tapbuf_L4SB_size8 mux_left_track_127 (
		.in({chany_bottom_in[62], left_bottom_grid_top_width_0_height_0_subtile_31__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_38__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_45__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_52__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_54__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_58__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_59__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_17_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_17_sram_inv[0:2]),
		.out(chanx_left_out[63]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_57 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size11_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_0_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_73 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size11_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_1_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_77 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size10_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_2_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_103 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size9_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_3_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_107 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size10_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_4_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_4_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_111 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size11_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_5_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_5_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_115 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size11_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_6_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_6_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_123 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size11_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_7_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_7_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_127 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size11_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_8_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_8_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_left_track_57 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size11_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_9_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_9_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_left_track_73 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size11_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_10_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_10_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_left_track_77 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size10_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_11_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_11_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_left_track_103 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size9_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_12_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_12_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_left_track_107 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size10_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_13_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_13_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_left_track_111 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size11_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_14_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_14_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_left_track_115 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size11_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_15_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_15_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_left_track_123 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size11_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_16_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_16_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_left_track_127 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size11_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_17_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_17_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size10 mux_bottom_track_75 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_27__pin_a2f_o_1_, chanx_left_in[38]}),
		.sram(mux_tree_tapbuf_L4SB_size10_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size10_0_sram_inv[0:3]),
		.out(chany_bottom_out[37]));

	mux_tree_tapbuf_L4SB_size10 mux_bottom_track_79 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_24__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_24__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_28__pin_a2f_o_1_, chanx_left_in[40]}),
		.sram(mux_tree_tapbuf_L4SB_size10_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size10_1_sram_inv[0:3]),
		.out(chany_bottom_out[39]));

	mux_tree_tapbuf_L4SB_size10 mux_bottom_track_83 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_25__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_25__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_29__pin_a2f_o_1_, chanx_left_in[42]}),
		.sram(mux_tree_tapbuf_L4SB_size10_2_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size10_2_sram_inv[0:3]),
		.out(chany_bottom_out[41]));

	mux_tree_tapbuf_L4SB_size10 mux_bottom_track_95 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_24__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_28__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_28__pin_a2f_o_1_, chanx_left_in[48]}),
		.sram(mux_tree_tapbuf_L4SB_size10_3_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size10_3_sram_inv[0:3]),
		.out(chany_bottom_out[47]));

	mux_tree_tapbuf_L4SB_size10 mux_bottom_track_99 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_25__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_29__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_29__pin_a2f_o_1_, chanx_left_in[50]}),
		.sram(mux_tree_tapbuf_L4SB_size10_4_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size10_4_sram_inv[0:3]),
		.out(chany_bottom_out[49]));

	mux_tree_tapbuf_L4SB_size10 mux_bottom_track_105 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_27__pin_a2f_o_0_, chanx_left_in[53]}),
		.sram(mux_tree_tapbuf_L4SB_size10_5_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size10_5_sram_inv[0:3]),
		.out(chany_bottom_out[52]));

	mux_tree_tapbuf_L4SB_size10 mux_bottom_track_117 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_, chanx_left_in[59]}),
		.sram(mux_tree_tapbuf_L4SB_size10_6_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size10_6_sram_inv[0:3]),
		.out(chany_bottom_out[58]));

	mux_tree_tapbuf_L4SB_size10 mux_left_track_75 (
		.in({chany_bottom_in[36], left_bottom_grid_top_width_0_height_0_subtile_32__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_39__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_41__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_45__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_46__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_49__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_53__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_53__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_57__pin_a2f_o_1_}),
		.sram(mux_tree_tapbuf_L4SB_size10_7_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size10_7_sram_inv[0:3]),
		.out(chanx_left_out[37]));

	mux_tree_tapbuf_L4SB_size10 mux_left_track_79 (
		.in({chany_bottom_in[38], left_bottom_grid_top_width_0_height_0_subtile_33__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_40__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_42__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_46__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_47__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_50__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_54__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_54__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_58__pin_a2f_o_1_}),
		.sram(mux_tree_tapbuf_L4SB_size10_8_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size10_8_sram_inv[0:3]),
		.out(chanx_left_out[39]));

	mux_tree_tapbuf_L4SB_size10 mux_left_track_83 (
		.in({chany_bottom_in[40], left_bottom_grid_top_width_0_height_0_subtile_34__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_41__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_43__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_47__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_48__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_51__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_55__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_55__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_59__pin_a2f_o_1_}),
		.sram(mux_tree_tapbuf_L4SB_size10_9_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size10_9_sram_inv[0:3]),
		.out(chanx_left_out[41]));

	mux_tree_tapbuf_L4SB_size10 mux_left_track_95 (
		.in({chany_bottom_in[46], left_bottom_grid_top_width_0_height_0_subtile_30__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_37__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_44__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_46__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_50__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_51__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_54__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_58__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_58__pin_a2f_o_1_}),
		.sram(mux_tree_tapbuf_L4SB_size10_10_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size10_10_sram_inv[0:3]),
		.out(chanx_left_out[47]));

	mux_tree_tapbuf_L4SB_size10 mux_left_track_99 (
		.in({chany_bottom_in[48], left_bottom_grid_top_width_0_height_0_subtile_31__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_38__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_45__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_47__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_51__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_52__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_55__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_59__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_59__pin_a2f_o_1_}),
		.sram(mux_tree_tapbuf_L4SB_size10_11_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size10_11_sram_inv[0:3]),
		.out(chanx_left_out[49]));

	mux_tree_tapbuf_L4SB_size10 mux_left_track_105 (
		.in({chany_bottom_in[51], left_bottom_grid_top_width_0_height_0_subtile_30__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_34__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_36__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_38__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_42__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_43__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_46__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_50__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_57__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size10_12_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size10_12_sram_inv[0:3]),
		.out(chanx_left_out[52]));

	mux_tree_tapbuf_L4SB_size10 mux_left_track_117 (
		.in({chany_bottom_in[57], left_bottom_grid_top_width_0_height_0_subtile_32__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_33__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_37__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_39__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_41__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_45__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_46__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_49__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_53__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size10_13_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size10_13_sram_inv[0:3]),
		.out(chanx_left_out[58]));

	mux_tree_tapbuf_L4SB_size10_mem mem_bottom_track_75 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size10_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size10_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size10_0_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size10_mem mem_bottom_track_79 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size10_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size10_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size10_1_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size10_mem mem_bottom_track_83 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size9_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size10_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size10_2_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size10_2_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size10_mem mem_bottom_track_95 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size9_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size10_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size10_3_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size10_3_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size10_mem mem_bottom_track_99 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size9_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size10_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size10_4_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size10_4_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size10_mem mem_bottom_track_105 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size10_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size10_5_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size10_5_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size10_mem mem_bottom_track_117 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size10_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size10_6_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size10_6_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size10_mem mem_left_track_75 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size10_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size10_7_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size10_7_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size10_mem mem_left_track_79 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size10_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size10_8_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size10_8_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size10_mem mem_left_track_83 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size9_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size10_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size10_9_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size10_9_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size10_mem mem_left_track_95 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size9_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size10_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size10_10_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size10_10_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size10_mem mem_left_track_99 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size9_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size10_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size10_11_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size10_11_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size10_mem mem_left_track_105 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size10_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size10_12_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size10_12_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size10_mem mem_left_track_117 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size10_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size10_13_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size10_13_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9 mux_bottom_track_81 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_21__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_28__pin_a2f_o_0_, chanx_left_in[41]}),
		.sram(mux_tree_tapbuf_L4SB_size9_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_0_sram_inv[0:3]),
		.out(chany_bottom_out[40]));

	mux_tree_tapbuf_L4SB_size9 mux_bottom_track_85 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_29__pin_a2f_o_0_, chanx_left_in[43]}),
		.sram(mux_tree_tapbuf_L4SB_size9_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_1_sram_inv[0:3]),
		.out(chany_bottom_out[42]));

	mux_tree_tapbuf_L4SB_size9 mux_bottom_track_87 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_26__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_26__pin_a2f_o_1_, chanx_left_in[44]}),
		.sram(mux_tree_tapbuf_L4SB_size9_2_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_2_sram_inv[0:3]),
		.out(chany_bottom_out[43]));

	mux_tree_tapbuf_L4SB_size9 mux_bottom_track_89 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_, chanx_left_in[45]}),
		.sram(mux_tree_tapbuf_L4SB_size9_3_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_3_sram_inv[0:3]),
		.out(chany_bottom_out[44]));

	mux_tree_tapbuf_L4SB_size9 mux_bottom_track_91 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_27__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_27__pin_a2f_o_1_, chanx_left_in[46]}),
		.sram(mux_tree_tapbuf_L4SB_size9_4_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_4_sram_inv[0:3]),
		.out(chany_bottom_out[45]));

	mux_tree_tapbuf_L4SB_size9 mux_bottom_track_93 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_24__pin_a2f_o_0_, chanx_left_in[47]}),
		.sram(mux_tree_tapbuf_L4SB_size9_5_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_5_sram_inv[0:3]),
		.out(chany_bottom_out[46]));

	mux_tree_tapbuf_L4SB_size9 mux_bottom_track_97 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_14__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_25__pin_a2f_o_0_, chanx_left_in[49]}),
		.sram(mux_tree_tapbuf_L4SB_size9_6_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_6_sram_inv[0:3]),
		.out(chany_bottom_out[48]));

	mux_tree_tapbuf_L4SB_size9 mux_bottom_track_101 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_26__pin_a2f_o_0_, chanx_left_in[51]}),
		.sram(mux_tree_tapbuf_L4SB_size9_7_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_7_sram_inv[0:3]),
		.out(chany_bottom_out[50]));

	mux_tree_tapbuf_L4SB_size9 mux_left_track_81 (
		.in({chany_bottom_in[39], left_bottom_grid_top_width_0_height_0_subtile_30__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_32__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_36__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_37__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_40__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_44__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_51__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_58__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size9_8_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_8_sram_inv[0:3]),
		.out(chanx_left_out[40]));

	mux_tree_tapbuf_L4SB_size9 mux_left_track_85 (
		.in({chany_bottom_in[41], left_bottom_grid_top_width_0_height_0_subtile_31__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_33__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_37__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_38__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_41__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_45__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_52__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_59__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size9_9_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_9_sram_inv[0:3]),
		.out(chanx_left_out[42]));

	mux_tree_tapbuf_L4SB_size9 mux_left_track_87 (
		.in({chany_bottom_in[42], left_bottom_grid_top_width_0_height_0_subtile_35__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_42__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_44__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_48__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_49__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_52__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_56__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_56__pin_a2f_o_1_}),
		.sram(mux_tree_tapbuf_L4SB_size9_10_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_10_sram_inv[0:3]),
		.out(chanx_left_out[43]));

	mux_tree_tapbuf_L4SB_size9 mux_left_track_89 (
		.in({chany_bottom_in[43], left_bottom_grid_top_width_0_height_0_subtile_30__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_32__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_34__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_38__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_39__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_42__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_46__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_53__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size9_11_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_11_sram_inv[0:3]),
		.out(chanx_left_out[44]));

	mux_tree_tapbuf_L4SB_size9 mux_left_track_91 (
		.in({chany_bottom_in[44], left_bottom_grid_top_width_0_height_0_subtile_36__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_43__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_45__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_49__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_50__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_53__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_57__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_57__pin_a2f_o_1_}),
		.sram(mux_tree_tapbuf_L4SB_size9_12_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_12_sram_inv[0:3]),
		.out(chanx_left_out[45]));

	mux_tree_tapbuf_L4SB_size9 mux_left_track_93 (
		.in({chany_bottom_in[45], left_bottom_grid_top_width_0_height_0_subtile_31__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_33__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_35__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_39__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_40__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_43__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_47__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_54__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size9_13_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_13_sram_inv[0:3]),
		.out(chanx_left_out[46]));

	mux_tree_tapbuf_L4SB_size9 mux_left_track_97 (
		.in({chany_bottom_in[47], left_bottom_grid_top_width_0_height_0_subtile_32__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_34__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_36__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_40__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_41__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_44__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_48__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_55__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size9_14_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_14_sram_inv[0:3]),
		.out(chanx_left_out[48]));

	mux_tree_tapbuf_L4SB_size9 mux_left_track_101 (
		.in({chany_bottom_in[49], left_bottom_grid_top_width_0_height_0_subtile_33__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_35__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_37__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_41__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_42__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_45__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_49__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_56__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size9_15_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size9_15_sram_inv[0:3]),
		.out(chanx_left_out[50]));

	mux_tree_tapbuf_L4SB_size9_mem mem_bottom_track_81 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size10_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size9_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size9_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_0_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_bottom_track_85 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size10_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size9_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size9_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_1_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_bottom_track_87 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size9_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size9_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size9_2_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_2_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_bottom_track_89 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size9_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size9_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size9_3_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_3_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_bottom_track_91 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size9_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size9_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size9_4_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_4_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_bottom_track_93 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size9_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size9_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size9_5_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_5_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_bottom_track_97 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size10_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size9_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size9_6_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_6_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_bottom_track_101 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size10_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size9_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size9_7_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_7_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_left_track_81 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size10_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size9_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size9_8_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_8_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_left_track_85 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size10_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size9_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size9_9_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_9_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_left_track_87 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size9_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size9_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size9_10_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_10_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_left_track_89 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size9_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size9_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size9_11_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_11_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_left_track_91 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size9_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size9_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size9_12_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_12_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_left_track_93 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size9_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size9_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size9_13_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_13_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_left_track_97 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size10_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size9_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size9_14_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_14_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size9_mem mem_left_track_101 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size10_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size9_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size9_15_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size9_15_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size5 mux_bottom_track_159 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_, chanx_left_in[80]}),
		.sram(mux_tree_tapbuf_L4SB_size5_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_0_sram_inv[0:2]),
		.out(chany_bottom_out[79]));

	mux_tree_tapbuf_L4SB_size5 mux_bottom_track_163 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_24__pin_a2f_o_0_, chanx_left_in[82]}),
		.sram(mux_tree_tapbuf_L4SB_size5_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_1_sram_inv[0:2]),
		.out(chany_bottom_out[81]));

	mux_tree_tapbuf_L4SB_size5 mux_bottom_track_167 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_11__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_18__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_25__pin_a2f_o_0_, chanx_left_in[84]}),
		.sram(mux_tree_tapbuf_L4SB_size5_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_2_sram_inv[0:2]),
		.out(chany_bottom_out[83]));

	mux_tree_tapbuf_L4SB_size5 mux_bottom_track_171 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_19__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_26__pin_a2f_o_0_, chanx_left_in[86]}),
		.sram(mux_tree_tapbuf_L4SB_size5_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_3_sram_inv[0:2]),
		.out(chany_bottom_out[85]));

	mux_tree_tapbuf_L4SB_size5 mux_bottom_track_175 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_13__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_27__pin_a2f_o_0_, chanx_left_in[88]}),
		.sram(mux_tree_tapbuf_L4SB_size5_4_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_4_sram_inv[0:2]),
		.out(chany_bottom_out[87]));

	mux_tree_tapbuf_L4SB_size5 mux_bottom_track_187 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_9__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_23__pin_a2f_o_0_, chanx_left_in[94]}),
		.sram(mux_tree_tapbuf_L4SB_size5_5_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_5_sram_inv[0:2]),
		.out(chany_bottom_out[93]));

	mux_tree_tapbuf_L4SB_size5 mux_bottom_track_191 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_10__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_17__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_24__pin_a2f_o_0_, chanx_left_in[0]}),
		.sram(mux_tree_tapbuf_L4SB_size5_6_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_6_sram_inv[0:2]),
		.out(chany_bottom_out[95]));

	mux_tree_tapbuf_L4SB_size5 mux_left_track_159 (
		.in({chany_bottom_in[78], left_bottom_grid_top_width_0_height_0_subtile_32__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_39__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_46__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_53__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size5_7_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_7_sram_inv[0:2]),
		.out(chanx_left_out[79]));

	mux_tree_tapbuf_L4SB_size5 mux_left_track_163 (
		.in({chany_bottom_in[80], left_bottom_grid_top_width_0_height_0_subtile_33__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_40__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_47__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_54__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size5_8_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_8_sram_inv[0:2]),
		.out(chanx_left_out[81]));

	mux_tree_tapbuf_L4SB_size5 mux_left_track_167 (
		.in({chany_bottom_in[82], left_bottom_grid_top_width_0_height_0_subtile_34__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_41__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_48__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_55__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size5_9_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_9_sram_inv[0:2]),
		.out(chanx_left_out[83]));

	mux_tree_tapbuf_L4SB_size5 mux_left_track_171 (
		.in({chany_bottom_in[84], left_bottom_grid_top_width_0_height_0_subtile_35__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_42__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_49__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_56__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size5_10_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_10_sram_inv[0:2]),
		.out(chanx_left_out[85]));

	mux_tree_tapbuf_L4SB_size5 mux_left_track_175 (
		.in({chany_bottom_in[86], left_bottom_grid_top_width_0_height_0_subtile_36__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_43__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_50__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_57__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size5_11_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_11_sram_inv[0:2]),
		.out(chanx_left_out[87]));

	mux_tree_tapbuf_L4SB_size5 mux_left_track_187 (
		.in({chany_bottom_in[92], left_bottom_grid_top_width_0_height_0_subtile_32__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_39__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_46__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_53__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size5_12_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_12_sram_inv[0:2]),
		.out(chanx_left_out[93]));

	mux_tree_tapbuf_L4SB_size5 mux_left_track_191 (
		.in({chany_bottom_in[94], left_bottom_grid_top_width_0_height_0_subtile_33__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_40__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_47__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_54__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size5_13_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size5_13_sram_inv[0:2]),
		.out(chanx_left_out[95]));

	mux_tree_tapbuf_L4SB_size5_mem mem_bottom_track_159 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size13_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size5_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size5_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_0_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size5_mem mem_bottom_track_163 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size12_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size5_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size5_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_1_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size5_mem mem_bottom_track_167 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size13_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size5_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size5_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_2_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size5_mem mem_bottom_track_171 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size14_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size5_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size5_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_3_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size5_mem mem_bottom_track_175 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size13_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size5_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size5_4_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_4_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size5_mem mem_bottom_track_187 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size13_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size5_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size5_5_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_5_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size5_mem mem_bottom_track_191 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size13_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size5_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size5_6_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_6_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size5_mem mem_left_track_159 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size13_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size5_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size5_7_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_7_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size5_mem mem_left_track_163 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size12_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size5_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size5_8_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_8_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size5_mem mem_left_track_167 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size13_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size5_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size5_9_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_9_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size5_mem mem_left_track_171 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size14_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size5_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size5_10_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_10_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size5_mem mem_left_track_175 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size13_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size5_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size5_11_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_11_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size5_mem mem_left_track_187 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size13_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size5_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size5_12_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_12_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size5_mem mem_left_track_191 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size13_mem_19_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size5_13_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size5_13_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size14 mux_bottom_track_169 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_8__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_12__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_15__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_16__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_20__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_22__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_24__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_28__pin_a2f_o_1_, bottom_left_grid_right_width_0_height_0_subtile_29__pin_a2f_o_0_, chanx_left_in[85]}),
		.sram(mux_tree_tapbuf_L4SB_size14_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size14_0_sram_inv[0:3]),
		.out(chany_bottom_out[84]));

	mux_tree_tapbuf_L4SB_size14 mux_left_track_169 (
		.in({chany_bottom_in[83], left_bottom_grid_top_width_0_height_0_subtile_30__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_31__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_34__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_38__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_38__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_42__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_45__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_46__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_50__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_52__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_54__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_58__pin_a2f_o_1_, left_bottom_grid_top_width_0_height_0_subtile_59__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size14_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_L4SB_size14_1_sram_inv[0:3]),
		.out(chanx_left_out[84]));

	mux_tree_tapbuf_L4SB_size14_mem mem_bottom_track_169 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size5_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size14_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size14_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size14_0_sram_inv[0:3]));

	mux_tree_tapbuf_L4SB_size14_mem mem_left_track_169 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size5_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size14_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size14_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_L4SB_size14_1_sram_inv[0:3]));

endmodule
// ----- END Verilog module for sb_10__8_ -----

//----- Default net type -----
`default_nettype none



