module add_1bit_1GE100_ES1(a, b, c);
input a, b;
output c;
                                 
  assign c = a + b;

endmodule  
