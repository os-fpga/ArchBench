//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for physical tile: bram]
//	Author: Xifan TANG
//	Organization: University of Utah
//-------------------------------------------
//----- Time scale -----
`timescale 1ns / 1ps

// ----- BEGIN Grid Verilog module: grid_bram -----
//----- Default net type -----
`default_nettype wire

// ----- Verilog module for grid_bram -----
module grid_bram(test_en,
                 scan_mode,
                 scan_clk,
                 config_enable,
                 prog_clock,
                 top_width_0_height_0_subtile_0__pin_PL_INIT_i_0_,
                 top_width_0_height_0_subtile_0__pin_PL_ENA_i_0_,
                 top_width_0_height_0_subtile_0__pin_PL_REN_i_0_,
                 top_width_0_height_0_subtile_0__pin_PL_WEN_i_0_,
                 top_width_0_height_0_subtile_0__pin_PL_WEN_i_1_,
                 top_width_0_height_0_subtile_0__pin_PL_ADDR_i_0_,
                 top_width_0_height_0_subtile_0__pin_PL_ADDR_i_1_,
                 top_width_0_height_0_subtile_0__pin_PL_ADDR_i_2_,
                 top_width_0_height_0_subtile_0__pin_PL_ADDR_i_3_,
                 top_width_0_height_0_subtile_0__pin_PL_ADDR_i_4_,
                 top_width_0_height_0_subtile_0__pin_PL_ADDR_i_5_,
                 top_width_0_height_0_subtile_0__pin_PL_ADDR_i_6_,
                 top_width_0_height_0_subtile_0__pin_PL_ADDR_i_7_,
                 top_width_0_height_0_subtile_0__pin_PL_ADDR_i_8_,
                 top_width_0_height_0_subtile_0__pin_PL_ADDR_i_9_,
                 top_width_0_height_0_subtile_0__pin_PL_ADDR_i_10_,
                 top_width_0_height_0_subtile_0__pin_PL_ADDR_i_11_,
                 top_width_0_height_0_subtile_0__pin_PL_ADDR_i_12_,
                 top_width_0_height_0_subtile_0__pin_PL_ADDR_i_13_,
                 top_width_0_height_0_subtile_0__pin_PL_ADDR_i_14_,
                 top_width_0_height_0_subtile_0__pin_PL_ADDR_i_15_,
                 top_width_0_height_0_subtile_0__pin_PL_ADDR_i_16_,
                 top_width_0_height_0_subtile_0__pin_PL_ADDR_i_17_,
                 top_width_0_height_0_subtile_0__pin_PL_ADDR_i_18_,
                 top_width_0_height_0_subtile_0__pin_PL_ADDR_i_19_,
                 top_width_0_height_0_subtile_0__pin_PL_ADDR_i_20_,
                 top_width_0_height_0_subtile_0__pin_PL_ADDR_i_21_,
                 top_width_0_height_0_subtile_0__pin_PL_ADDR_i_22_,
                 top_width_0_height_0_subtile_0__pin_PL_ADDR_i_23_,
                 top_width_0_height_0_subtile_0__pin_PL_ADDR_i_24_,
                 top_width_0_height_0_subtile_0__pin_PL_ADDR_i_25_,
                 top_width_0_height_0_subtile_0__pin_PL_ADDR_i_26_,
                 top_width_0_height_0_subtile_0__pin_PL_ADDR_i_27_,
                 top_width_0_height_0_subtile_0__pin_PL_ADDR_i_28_,
                 top_width_0_height_0_subtile_0__pin_PL_ADDR_i_29_,
                 top_width_0_height_0_subtile_0__pin_PL_ADDR_i_30_,
                 top_width_0_height_0_subtile_0__pin_PL_ADDR_i_31_,
                 top_width_0_height_0_subtile_0__pin_PL_DATA_i_0_,
                 top_width_0_height_0_subtile_0__pin_PL_DATA_i_1_,
                 top_width_0_height_0_subtile_0__pin_PL_DATA_i_2_,
                 top_width_0_height_0_subtile_0__pin_PL_DATA_i_3_,
                 top_width_0_height_0_subtile_0__pin_PL_DATA_i_4_,
                 top_width_0_height_0_subtile_0__pin_PL_DATA_i_5_,
                 top_width_0_height_0_subtile_0__pin_PL_DATA_i_6_,
                 top_width_0_height_0_subtile_0__pin_PL_DATA_i_7_,
                 top_width_0_height_0_subtile_0__pin_PL_DATA_i_8_,
                 top_width_0_height_0_subtile_0__pin_PL_DATA_i_9_,
                 top_width_0_height_0_subtile_0__pin_PL_DATA_i_10_,
                 top_width_0_height_0_subtile_0__pin_PL_DATA_i_11_,
                 top_width_0_height_0_subtile_0__pin_PL_DATA_i_12_,
                 top_width_0_height_0_subtile_0__pin_PL_DATA_i_13_,
                 top_width_0_height_0_subtile_0__pin_PL_DATA_i_14_,
                 top_width_0_height_0_subtile_0__pin_PL_DATA_i_15_,
                 top_width_0_height_0_subtile_0__pin_PL_DATA_i_16_,
                 top_width_0_height_0_subtile_0__pin_PL_DATA_i_17_,
                 top_width_0_height_0_subtile_0__pin_PL_DATA_i_18_,
                 top_width_0_height_0_subtile_0__pin_PL_DATA_i_19_,
                 top_width_0_height_0_subtile_0__pin_PL_DATA_i_20_,
                 top_width_0_height_0_subtile_0__pin_PL_DATA_i_21_,
                 top_width_0_height_0_subtile_0__pin_PL_DATA_i_22_,
                 top_width_0_height_0_subtile_0__pin_PL_DATA_i_23_,
                 top_width_0_height_0_subtile_0__pin_PL_DATA_i_24_,
                 top_width_0_height_0_subtile_0__pin_PL_DATA_i_25_,
                 top_width_0_height_0_subtile_0__pin_PL_DATA_i_26_,
                 top_width_0_height_0_subtile_0__pin_PL_DATA_i_27_,
                 top_width_0_height_0_subtile_0__pin_PL_DATA_i_28_,
                 top_width_0_height_0_subtile_0__pin_PL_DATA_i_29_,
                 top_width_0_height_0_subtile_0__pin_PL_DATA_i_30_,
                 top_width_0_height_0_subtile_0__pin_PL_DATA_i_31_,
                 top_width_0_height_0_subtile_0__pin_PL_DATA_i_32_,
                 top_width_0_height_0_subtile_0__pin_PL_DATA_i_33_,
                 top_width_0_height_0_subtile_0__pin_PL_DATA_i_34_,
                 top_width_0_height_0_subtile_0__pin_PL_DATA_i_35_,
                 top_width_0_height_0_subtile_0__pin_sc_in_0_,
                 top_width_0_height_0_subtile_0__pin_sc_in_1_,
                 top_width_0_height_0_subtile_0__pin_sc_in_2_,
                 top_width_0_height_0_subtile_0__pin_sc_in_3_,
                 top_width_0_height_0_subtile_0__pin_sc_in_4_,
                 top_width_0_height_0_subtile_0__pin_sc_in_5_,
                 top_width_0_height_0_subtile_0__pin_PL_CLK_i_0_,
                 right_width_0_height_0_subtile_0__pin_ADDR_A1_i_2_,
                 right_width_0_height_0_subtile_0__pin_ADDR_A1_i_3_,
                 right_width_0_height_0_subtile_0__pin_ADDR_A1_i_4_,
                 right_width_0_height_0_subtile_0__pin_ADDR_A1_i_5_,
                 right_width_0_height_0_subtile_0__pin_WDATA_B1_i_1_,
                 right_width_0_height_0_subtile_0__pin_WDATA_B1_i_2_,
                 right_width_0_height_0_subtile_0__pin_WDATA_B1_i_3_,
                 right_width_0_height_0_subtile_0__pin_WDATA_B1_i_4_,
                 right_width_0_height_0_subtile_0__pin_WDATA_B1_i_5_,
                 right_width_0_height_0_subtile_0__pin_WDATA_B1_i_6_,
                 right_width_0_height_0_subtile_0__pin_WDATA_B1_i_7_,
                 right_width_0_height_0_subtile_0__pin_WDATA_B1_i_8_,
                 right_width_0_height_0_subtile_0__pin_WDATA_B1_i_9_,
                 right_width_0_height_0_subtile_0__pin_WDATA_B1_i_10_,
                 right_width_0_height_0_subtile_0__pin_WDATA_B1_i_11_,
                 right_width_0_height_0_subtile_0__pin_WDATA_B1_i_12_,
                 right_width_0_height_0_subtile_0__pin_WDATA_B1_i_13_,
                 right_width_0_height_0_subtile_0__pin_WDATA_B1_i_14_,
                 right_width_0_height_0_subtile_0__pin_WDATA_B1_i_15_,
                 right_width_0_height_0_subtile_0__pin_WDATA_B1_i_16_,
                 right_width_0_height_0_subtile_0__pin_ADDR_B1_i_0_,
                 right_width_0_height_1_subtile_0__pin_WDATA_A2_i_17_,
                 right_width_0_height_1_subtile_0__pin_ADDR_A2_i_1_,
                 right_width_0_height_1_subtile_0__pin_REN_A1_i_0_,
                 right_width_0_height_1_subtile_0__pin_REN_A2_i_0_,
                 right_width_0_height_1_subtile_0__pin_WEN_A2_i_0_,
                 right_width_0_height_1_subtile_0__pin_BE_A2_i_0_,
                 right_width_0_height_1_subtile_0__pin_BE_A2_i_1_,
                 right_width_0_height_1_subtile_0__pin_WDATA_B1_i_0_,
                 right_width_0_height_1_subtile_0__pin_ADDR_B1_i_2_,
                 right_width_0_height_1_subtile_0__pin_ADDR_B1_i_3_,
                 right_width_0_height_1_subtile_0__pin_ADDR_B1_i_4_,
                 right_width_0_height_1_subtile_0__pin_ADDR_B1_i_5_,
                 right_width_0_height_1_subtile_0__pin_ADDR_B1_i_6_,
                 right_width_0_height_1_subtile_0__pin_ADDR_B1_i_7_,
                 right_width_0_height_1_subtile_0__pin_ADDR_B1_i_8_,
                 right_width_0_height_1_subtile_0__pin_ADDR_B1_i_9_,
                 right_width_0_height_1_subtile_0__pin_ADDR_B1_i_10_,
                 right_width_0_height_1_subtile_0__pin_ADDR_B1_i_11_,
                 right_width_0_height_1_subtile_0__pin_ADDR_B1_i_12_,
                 right_width_0_height_1_subtile_0__pin_ADDR_B1_i_13_,
                 right_width_0_height_1_subtile_0__pin_ADDR_B1_i_14_,
                 right_width_0_height_1_subtile_0__pin_FLUSH2_i_0_,
                 right_width_0_height_2_subtile_0__pin_WDATA_A2_i_9_,
                 right_width_0_height_2_subtile_0__pin_WDATA_A2_i_10_,
                 right_width_0_height_2_subtile_0__pin_WDATA_A2_i_11_,
                 right_width_0_height_2_subtile_0__pin_WDATA_A2_i_12_,
                 right_width_0_height_2_subtile_0__pin_WDATA_A2_i_13_,
                 right_width_0_height_2_subtile_0__pin_WDATA_A2_i_14_,
                 right_width_0_height_2_subtile_0__pin_WDATA_A2_i_15_,
                 right_width_0_height_2_subtile_0__pin_WDATA_A2_i_16_,
                 right_width_0_height_2_subtile_0__pin_ADDR_A2_i_0_,
                 right_width_0_height_2_subtile_0__pin_ADDR_A2_i_2_,
                 right_width_0_height_2_subtile_0__pin_ADDR_A2_i_3_,
                 right_width_0_height_2_subtile_0__pin_ADDR_A2_i_4_,
                 right_width_0_height_2_subtile_0__pin_ADDR_A2_i_5_,
                 right_width_0_height_2_subtile_0__pin_ADDR_A2_i_6_,
                 right_width_0_height_2_subtile_0__pin_ADDR_A2_i_7_,
                 right_width_0_height_2_subtile_0__pin_ADDR_A2_i_8_,
                 right_width_0_height_2_subtile_0__pin_ADDR_A2_i_9_,
                 right_width_0_height_2_subtile_0__pin_ADDR_A2_i_10_,
                 right_width_0_height_2_subtile_0__pin_ADDR_A2_i_11_,
                 right_width_0_height_2_subtile_0__pin_ADDR_A2_i_12_,
                 right_width_0_height_2_subtile_0__pin_ADDR_A2_i_13_,
                 right_width_0_height_2_subtile_0__pin_WEN_A1_i_0_,
                 right_width_0_height_3_subtile_0__pin_WDATA_A1_i_7_,
                 right_width_0_height_3_subtile_0__pin_WDATA_A1_i_8_,
                 right_width_0_height_3_subtile_0__pin_WDATA_A1_i_9_,
                 right_width_0_height_3_subtile_0__pin_WDATA_A1_i_10_,
                 right_width_0_height_3_subtile_0__pin_WDATA_A1_i_11_,
                 right_width_0_height_3_subtile_0__pin_WDATA_A1_i_12_,
                 right_width_0_height_3_subtile_0__pin_WDATA_A1_i_13_,
                 right_width_0_height_3_subtile_0__pin_WDATA_A1_i_14_,
                 right_width_0_height_3_subtile_0__pin_WDATA_A1_i_15_,
                 right_width_0_height_3_subtile_0__pin_WDATA_A1_i_16_,
                 right_width_0_height_3_subtile_0__pin_WDATA_A1_i_17_,
                 right_width_0_height_3_subtile_0__pin_ADDR_A1_i_0_,
                 right_width_0_height_3_subtile_0__pin_ADDR_A1_i_1_,
                 right_width_0_height_3_subtile_0__pin_BE_A1_i_0_,
                 right_width_0_height_3_subtile_0__pin_BE_A1_i_1_,
                 right_width_0_height_3_subtile_0__pin_REN_B2_i_0_,
                 right_width_0_height_3_subtile_0__pin_WEN_B2_i_0_,
                 right_width_0_height_3_subtile_0__pin_BE_B1_i_0_,
                 right_width_0_height_3_subtile_0__pin_BE_B1_i_1_,
                 right_width_0_height_3_subtile_0__pin_BE_B2_i_0_,
                 right_width_0_height_3_subtile_0__pin_BE_B2_i_1_,
                 right_width_0_height_3_subtile_0__pin_FLUSH1_i_0_,
                 right_width_0_height_4_subtile_0__pin_WDATA_A2_i_0_,
                 right_width_0_height_4_subtile_0__pin_WDATA_A2_i_1_,
                 right_width_0_height_4_subtile_0__pin_WDATA_A2_i_2_,
                 right_width_0_height_4_subtile_0__pin_WDATA_A2_i_3_,
                 right_width_0_height_4_subtile_0__pin_WDATA_A2_i_4_,
                 right_width_0_height_4_subtile_0__pin_WDATA_A2_i_5_,
                 right_width_0_height_4_subtile_0__pin_WDATA_A2_i_6_,
                 right_width_0_height_4_subtile_0__pin_WDATA_A2_i_7_,
                 right_width_0_height_4_subtile_0__pin_WDATA_A2_i_8_,
                 right_width_0_height_4_subtile_0__pin_WDATA_B2_i_17_,
                 right_width_0_height_4_subtile_0__pin_ADDR_B2_i_1_,
                 right_width_0_height_4_subtile_0__pin_ADDR_B2_i_4_,
                 right_width_0_height_4_subtile_0__pin_ADDR_B2_i_5_,
                 right_width_0_height_4_subtile_0__pin_ADDR_B2_i_6_,
                 right_width_0_height_4_subtile_0__pin_ADDR_B2_i_7_,
                 right_width_0_height_4_subtile_0__pin_ADDR_B2_i_8_,
                 right_width_0_height_4_subtile_0__pin_ADDR_B2_i_9_,
                 right_width_0_height_4_subtile_0__pin_ADDR_B2_i_10_,
                 right_width_0_height_4_subtile_0__pin_ADDR_B2_i_11_,
                 right_width_0_height_4_subtile_0__pin_ADDR_B2_i_12_,
                 right_width_0_height_4_subtile_0__pin_ADDR_B2_i_13_,
                 right_width_0_height_4_subtile_0__pin_WEN_B1_i_0_,
                 right_width_0_height_5_subtile_0__pin_WDATA_B2_i_0_,
                 right_width_0_height_5_subtile_0__pin_WDATA_B2_i_1_,
                 right_width_0_height_5_subtile_0__pin_WDATA_B2_i_2_,
                 right_width_0_height_5_subtile_0__pin_WDATA_B2_i_3_,
                 right_width_0_height_5_subtile_0__pin_WDATA_B2_i_4_,
                 right_width_0_height_5_subtile_0__pin_WDATA_B2_i_5_,
                 right_width_0_height_5_subtile_0__pin_WDATA_B2_i_6_,
                 right_width_0_height_5_subtile_0__pin_WDATA_B2_i_7_,
                 right_width_0_height_5_subtile_0__pin_WDATA_B2_i_8_,
                 right_width_0_height_5_subtile_0__pin_WDATA_B2_i_9_,
                 right_width_0_height_5_subtile_0__pin_WDATA_B2_i_10_,
                 right_width_0_height_5_subtile_0__pin_WDATA_B2_i_11_,
                 right_width_0_height_5_subtile_0__pin_WDATA_B2_i_12_,
                 right_width_0_height_5_subtile_0__pin_WDATA_B2_i_13_,
                 right_width_0_height_5_subtile_0__pin_WDATA_B2_i_14_,
                 right_width_0_height_5_subtile_0__pin_WDATA_B2_i_15_,
                 right_width_0_height_5_subtile_0__pin_WDATA_B2_i_16_,
                 right_width_0_height_5_subtile_0__pin_ADDR_B2_i_0_,
                 right_width_0_height_5_subtile_0__pin_ADDR_B2_i_2_,
                 right_width_0_height_5_subtile_0__pin_ADDR_B2_i_3_,
                 right_width_0_height_5_subtile_0__pin_REN_B1_i_0_,
                 bottom_width_0_height_0_subtile_0__pin_WDATA_A1_i_0_,
                 bottom_width_0_height_0_subtile_0__pin_WDATA_A1_i_1_,
                 bottom_width_0_height_0_subtile_0__pin_WDATA_A1_i_2_,
                 bottom_width_0_height_0_subtile_0__pin_WDATA_A1_i_3_,
                 bottom_width_0_height_0_subtile_0__pin_WDATA_A1_i_4_,
                 bottom_width_0_height_0_subtile_0__pin_WDATA_A1_i_5_,
                 bottom_width_0_height_0_subtile_0__pin_WDATA_A1_i_6_,
                 bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_6_,
                 bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_7_,
                 bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_8_,
                 bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_9_,
                 bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_10_,
                 bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_11_,
                 bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_12_,
                 bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_13_,
                 bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_14_,
                 bottom_width_0_height_0_subtile_0__pin_WDATA_B1_i_17_,
                 bottom_width_0_height_0_subtile_0__pin_ADDR_B1_i_1_,
                 left_width_0_height_0_subtile_0__pin_RAM_ID_i_0_,
                 left_width_0_height_0_subtile_0__pin_RAM_ID_i_1_,
                 left_width_0_height_0_subtile_0__pin_RAM_ID_i_2_,
                 left_width_0_height_0_subtile_0__pin_RAM_ID_i_3_,
                 left_width_0_height_0_subtile_0__pin_RAM_ID_i_4_,
                 left_width_0_height_0_subtile_0__pin_RAM_ID_i_5_,
                 left_width_0_height_0_subtile_0__pin_RAM_ID_i_6_,
                 left_width_0_height_0_subtile_0__pin_RAM_ID_i_7_,
                 left_width_0_height_0_subtile_0__pin_RAM_ID_i_8_,
                 left_width_0_height_0_subtile_0__pin_RAM_ID_i_9_,
                 left_width_0_height_0_subtile_0__pin_RAM_ID_i_10_,
                 left_width_0_height_0_subtile_0__pin_RAM_ID_i_11_,
                 left_width_0_height_0_subtile_0__pin_RAM_ID_i_12_,
                 left_width_0_height_0_subtile_0__pin_RAM_ID_i_13_,
                 left_width_0_height_0_subtile_0__pin_RAM_ID_i_14_,
                 left_width_0_height_0_subtile_0__pin_RAM_ID_i_15_,
                 left_width_0_height_0_subtile_0__pin_RAM_ID_i_16_,
                 left_width_0_height_0_subtile_0__pin_RAM_ID_i_17_,
                 left_width_0_height_0_subtile_0__pin_RAM_ID_i_18_,
                 left_width_0_height_0_subtile_0__pin_RAM_ID_i_19_,
                 left_width_0_height_0_subtile_0__pin_global_reset_0_,
                 left_width_0_height_0_subtile_0__pin_scan_reset_0_,
                 left_width_0_height_0_subtile_0__pin_clk_0_,
                 left_width_0_height_0_subtile_0__pin_clk_1_,
                 left_width_0_height_0_subtile_0__pin_clk_2_,
                 left_width_0_height_0_subtile_0__pin_clk_3_,
                 ccff_head,
                 right_width_0_height_0_subtile_0__pin_RDATA_A1_o_0_,
                 right_width_0_height_0_subtile_0__pin_RDATA_A1_o_1_,
                 right_width_0_height_0_subtile_0__pin_RDATA_A1_o_2_,
                 right_width_0_height_0_subtile_0__pin_RDATA_A1_o_3_,
                 right_width_0_height_0_subtile_0__pin_RDATA_A1_o_4_,
                 right_width_0_height_0_subtile_0__pin_RDATA_A1_o_5_,
                 right_width_0_height_0_subtile_0__pin_RDATA_B1_o_0_,
                 right_width_0_height_0_subtile_0__pin_RDATA_B1_o_1_,
                 right_width_0_height_0_subtile_0__pin_RDATA_B1_o_2_,
                 right_width_0_height_0_subtile_0__pin_RDATA_B1_o_3_,
                 right_width_0_height_0_subtile_0__pin_RDATA_B1_o_4_,
                 right_width_0_height_0_subtile_0__pin_RDATA_B1_o_5_,
                 right_width_0_height_1_subtile_0__pin_RDATA_A1_o_6_,
                 right_width_0_height_1_subtile_0__pin_RDATA_A1_o_7_,
                 right_width_0_height_1_subtile_0__pin_RDATA_A1_o_8_,
                 right_width_0_height_1_subtile_0__pin_RDATA_A1_o_9_,
                 right_width_0_height_1_subtile_0__pin_RDATA_A1_o_10_,
                 right_width_0_height_1_subtile_0__pin_RDATA_A1_o_11_,
                 right_width_0_height_1_subtile_0__pin_RDATA_B1_o_6_,
                 right_width_0_height_1_subtile_0__pin_RDATA_B1_o_7_,
                 right_width_0_height_1_subtile_0__pin_RDATA_B1_o_8_,
                 right_width_0_height_1_subtile_0__pin_RDATA_B1_o_9_,
                 right_width_0_height_1_subtile_0__pin_RDATA_B1_o_10_,
                 right_width_0_height_1_subtile_0__pin_RDATA_B1_o_11_,
                 right_width_0_height_2_subtile_0__pin_RDATA_A1_o_12_,
                 right_width_0_height_2_subtile_0__pin_RDATA_A1_o_13_,
                 right_width_0_height_2_subtile_0__pin_RDATA_A1_o_14_,
                 right_width_0_height_2_subtile_0__pin_RDATA_A1_o_15_,
                 right_width_0_height_2_subtile_0__pin_RDATA_A1_o_16_,
                 right_width_0_height_2_subtile_0__pin_RDATA_A1_o_17_,
                 right_width_0_height_2_subtile_0__pin_RDATA_B1_o_12_,
                 right_width_0_height_2_subtile_0__pin_RDATA_B1_o_13_,
                 right_width_0_height_2_subtile_0__pin_RDATA_B1_o_14_,
                 right_width_0_height_2_subtile_0__pin_RDATA_B1_o_15_,
                 right_width_0_height_2_subtile_0__pin_RDATA_B1_o_16_,
                 right_width_0_height_2_subtile_0__pin_RDATA_B1_o_17_,
                 right_width_0_height_3_subtile_0__pin_RDATA_A2_o_0_,
                 right_width_0_height_3_subtile_0__pin_RDATA_A2_o_1_,
                 right_width_0_height_3_subtile_0__pin_RDATA_A2_o_2_,
                 right_width_0_height_3_subtile_0__pin_RDATA_A2_o_3_,
                 right_width_0_height_3_subtile_0__pin_RDATA_A2_o_4_,
                 right_width_0_height_3_subtile_0__pin_RDATA_A2_o_5_,
                 right_width_0_height_3_subtile_0__pin_RDATA_B2_o_0_,
                 right_width_0_height_3_subtile_0__pin_RDATA_B2_o_1_,
                 right_width_0_height_3_subtile_0__pin_RDATA_B2_o_2_,
                 right_width_0_height_3_subtile_0__pin_RDATA_B2_o_3_,
                 right_width_0_height_3_subtile_0__pin_RDATA_B2_o_4_,
                 right_width_0_height_3_subtile_0__pin_RDATA_B2_o_5_,
                 right_width_0_height_4_subtile_0__pin_RDATA_A2_o_6_,
                 right_width_0_height_4_subtile_0__pin_RDATA_A2_o_7_,
                 right_width_0_height_4_subtile_0__pin_RDATA_A2_o_8_,
                 right_width_0_height_4_subtile_0__pin_RDATA_A2_o_9_,
                 right_width_0_height_4_subtile_0__pin_RDATA_A2_o_10_,
                 right_width_0_height_4_subtile_0__pin_RDATA_A2_o_11_,
                 right_width_0_height_4_subtile_0__pin_RDATA_B2_o_6_,
                 right_width_0_height_4_subtile_0__pin_RDATA_B2_o_7_,
                 right_width_0_height_4_subtile_0__pin_RDATA_B2_o_8_,
                 right_width_0_height_4_subtile_0__pin_RDATA_B2_o_9_,
                 right_width_0_height_4_subtile_0__pin_RDATA_B2_o_10_,
                 right_width_0_height_4_subtile_0__pin_RDATA_B2_o_11_,
                 right_width_0_height_5_subtile_0__pin_RDATA_A2_o_12_,
                 right_width_0_height_5_subtile_0__pin_RDATA_A2_o_13_,
                 right_width_0_height_5_subtile_0__pin_RDATA_A2_o_14_,
                 right_width_0_height_5_subtile_0__pin_RDATA_A2_o_15_,
                 right_width_0_height_5_subtile_0__pin_RDATA_A2_o_16_,
                 right_width_0_height_5_subtile_0__pin_RDATA_A2_o_17_,
                 right_width_0_height_5_subtile_0__pin_RDATA_B2_o_12_,
                 right_width_0_height_5_subtile_0__pin_RDATA_B2_o_13_,
                 right_width_0_height_5_subtile_0__pin_RDATA_B2_o_14_,
                 right_width_0_height_5_subtile_0__pin_RDATA_B2_o_15_,
                 right_width_0_height_5_subtile_0__pin_RDATA_B2_o_16_,
                 right_width_0_height_5_subtile_0__pin_RDATA_B2_o_17_,
                 bottom_width_0_height_0_subtile_0__pin_PL_INIT_o_0_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ENA_o_0_,
                 bottom_width_0_height_0_subtile_0__pin_PL_REN_o_0_,
                 bottom_width_0_height_0_subtile_0__pin_PL_CLK_o_0_,
                 bottom_width_0_height_0_subtile_0__pin_PL_WEN_o_0_,
                 bottom_width_0_height_0_subtile_0__pin_PL_WEN_o_1_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_0_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_1_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_2_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_3_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_4_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_5_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_6_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_7_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_8_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_9_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_10_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_11_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_12_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_13_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_14_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_15_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_16_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_17_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_18_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_19_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_20_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_21_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_22_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_23_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_24_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_25_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_26_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_27_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_28_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_29_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_30_,
                 bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_31_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_0_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_1_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_2_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_3_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_4_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_5_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_6_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_7_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_8_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_9_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_10_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_11_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_12_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_13_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_14_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_15_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_16_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_17_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_18_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_19_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_20_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_21_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_22_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_23_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_24_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_25_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_26_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_27_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_28_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_29_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_30_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_31_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_32_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_33_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_34_,
                 bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_35_,
                 bottom_width_0_height_0_subtile_0__pin_sc_out_0_,
                 bottom_width_0_height_0_subtile_0__pin_sc_out_1_,
                 bottom_width_0_height_0_subtile_0__pin_sc_out_2_,
                 bottom_width_0_height_0_subtile_0__pin_sc_out_3_,
                 bottom_width_0_height_0_subtile_0__pin_sc_out_4_,
                 bottom_width_0_height_0_subtile_0__pin_sc_out_5_,
                 ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] test_en;
//----- GLOBAL PORTS -----
input [0:0] scan_mode;
//----- GLOBAL PORTS -----
input [0:0] scan_clk;
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_clock;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_INIT_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_ENA_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_REN_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_WEN_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_WEN_i_1_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_ADDR_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_ADDR_i_1_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_ADDR_i_2_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_ADDR_i_3_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_ADDR_i_4_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_ADDR_i_5_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_ADDR_i_6_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_ADDR_i_7_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_ADDR_i_8_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_ADDR_i_9_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_ADDR_i_10_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_ADDR_i_11_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_ADDR_i_12_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_ADDR_i_13_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_ADDR_i_14_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_ADDR_i_15_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_ADDR_i_16_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_ADDR_i_17_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_ADDR_i_18_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_ADDR_i_19_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_ADDR_i_20_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_ADDR_i_21_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_ADDR_i_22_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_ADDR_i_23_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_ADDR_i_24_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_ADDR_i_25_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_ADDR_i_26_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_ADDR_i_27_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_ADDR_i_28_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_ADDR_i_29_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_ADDR_i_30_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_ADDR_i_31_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_DATA_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_DATA_i_1_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_DATA_i_2_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_DATA_i_3_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_DATA_i_4_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_DATA_i_5_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_DATA_i_6_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_DATA_i_7_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_DATA_i_8_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_DATA_i_9_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_DATA_i_10_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_DATA_i_11_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_DATA_i_12_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_DATA_i_13_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_DATA_i_14_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_DATA_i_15_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_DATA_i_16_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_DATA_i_17_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_DATA_i_18_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_DATA_i_19_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_DATA_i_20_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_DATA_i_21_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_DATA_i_22_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_DATA_i_23_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_DATA_i_24_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_DATA_i_25_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_DATA_i_26_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_DATA_i_27_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_DATA_i_28_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_DATA_i_29_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_DATA_i_30_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_DATA_i_31_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_DATA_i_32_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_DATA_i_33_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_DATA_i_34_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_DATA_i_35_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_sc_in_1_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_sc_in_2_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_sc_in_3_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_sc_in_4_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_sc_in_5_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_PL_CLK_i_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_ADDR_A1_i_2_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_ADDR_A1_i_3_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_ADDR_A1_i_4_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_ADDR_A1_i_5_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_WDATA_B1_i_1_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_WDATA_B1_i_2_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_WDATA_B1_i_3_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_WDATA_B1_i_4_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_WDATA_B1_i_5_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_WDATA_B1_i_6_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_WDATA_B1_i_7_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_WDATA_B1_i_8_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_WDATA_B1_i_9_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_WDATA_B1_i_10_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_WDATA_B1_i_11_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_WDATA_B1_i_12_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_WDATA_B1_i_13_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_WDATA_B1_i_14_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_WDATA_B1_i_15_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_WDATA_B1_i_16_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_ADDR_B1_i_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_WDATA_A2_i_17_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_ADDR_A2_i_1_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_REN_A1_i_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_REN_A2_i_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_WEN_A2_i_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_BE_A2_i_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_BE_A2_i_1_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_WDATA_B1_i_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_ADDR_B1_i_2_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_ADDR_B1_i_3_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_ADDR_B1_i_4_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_ADDR_B1_i_5_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_ADDR_B1_i_6_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_ADDR_B1_i_7_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_ADDR_B1_i_8_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_ADDR_B1_i_9_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_ADDR_B1_i_10_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_ADDR_B1_i_11_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_ADDR_B1_i_12_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_ADDR_B1_i_13_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_ADDR_B1_i_14_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_1_subtile_0__pin_FLUSH2_i_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_WDATA_A2_i_9_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_WDATA_A2_i_10_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_WDATA_A2_i_11_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_WDATA_A2_i_12_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_WDATA_A2_i_13_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_WDATA_A2_i_14_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_WDATA_A2_i_15_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_WDATA_A2_i_16_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_ADDR_A2_i_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_ADDR_A2_i_2_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_ADDR_A2_i_3_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_ADDR_A2_i_4_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_ADDR_A2_i_5_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_ADDR_A2_i_6_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_ADDR_A2_i_7_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_ADDR_A2_i_8_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_ADDR_A2_i_9_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_ADDR_A2_i_10_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_ADDR_A2_i_11_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_ADDR_A2_i_12_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_ADDR_A2_i_13_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_2_subtile_0__pin_WEN_A1_i_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_WDATA_A1_i_7_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_WDATA_A1_i_8_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_WDATA_A1_i_9_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_WDATA_A1_i_10_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_WDATA_A1_i_11_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_WDATA_A1_i_12_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_WDATA_A1_i_13_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_WDATA_A1_i_14_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_WDATA_A1_i_15_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_WDATA_A1_i_16_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_WDATA_A1_i_17_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_ADDR_A1_i_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_ADDR_A1_i_1_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_BE_A1_i_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_BE_A1_i_1_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_REN_B2_i_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_WEN_B2_i_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_BE_B1_i_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_BE_B1_i_1_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_BE_B2_i_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_BE_B2_i_1_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_3_subtile_0__pin_FLUSH1_i_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_4_subtile_0__pin_WDATA_A2_i_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_4_subtile_0__pin_WDATA_A2_i_1_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_4_subtile_0__pin_WDATA_A2_i_2_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_4_subtile_0__pin_WDATA_A2_i_3_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_4_subtile_0__pin_WDATA_A2_i_4_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_4_subtile_0__pin_WDATA_A2_i_5_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_4_subtile_0__pin_WDATA_A2_i_6_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_4_subtile_0__pin_WDATA_A2_i_7_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_4_subtile_0__pin_WDATA_A2_i_8_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_4_subtile_0__pin_WDATA_B2_i_17_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_4_subtile_0__pin_ADDR_B2_i_1_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_4_subtile_0__pin_ADDR_B2_i_4_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_4_subtile_0__pin_ADDR_B2_i_5_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_4_subtile_0__pin_ADDR_B2_i_6_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_4_subtile_0__pin_ADDR_B2_i_7_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_4_subtile_0__pin_ADDR_B2_i_8_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_4_subtile_0__pin_ADDR_B2_i_9_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_4_subtile_0__pin_ADDR_B2_i_10_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_4_subtile_0__pin_ADDR_B2_i_11_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_4_subtile_0__pin_ADDR_B2_i_12_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_4_subtile_0__pin_ADDR_B2_i_13_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_4_subtile_0__pin_WEN_B1_i_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_5_subtile_0__pin_WDATA_B2_i_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_5_subtile_0__pin_WDATA_B2_i_1_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_5_subtile_0__pin_WDATA_B2_i_2_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_5_subtile_0__pin_WDATA_B2_i_3_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_5_subtile_0__pin_WDATA_B2_i_4_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_5_subtile_0__pin_WDATA_B2_i_5_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_5_subtile_0__pin_WDATA_B2_i_6_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_5_subtile_0__pin_WDATA_B2_i_7_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_5_subtile_0__pin_WDATA_B2_i_8_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_5_subtile_0__pin_WDATA_B2_i_9_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_5_subtile_0__pin_WDATA_B2_i_10_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_5_subtile_0__pin_WDATA_B2_i_11_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_5_subtile_0__pin_WDATA_B2_i_12_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_5_subtile_0__pin_WDATA_B2_i_13_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_5_subtile_0__pin_WDATA_B2_i_14_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_5_subtile_0__pin_WDATA_B2_i_15_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_5_subtile_0__pin_WDATA_B2_i_16_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_5_subtile_0__pin_ADDR_B2_i_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_5_subtile_0__pin_ADDR_B2_i_2_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_5_subtile_0__pin_ADDR_B2_i_3_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_5_subtile_0__pin_REN_B1_i_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_WDATA_A1_i_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_WDATA_A1_i_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_WDATA_A1_i_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_WDATA_A1_i_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_WDATA_A1_i_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_WDATA_A1_i_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_WDATA_A1_i_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_WDATA_B1_i_17_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_ADDR_B1_i_1_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_RAM_ID_i_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_RAM_ID_i_1_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_RAM_ID_i_2_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_RAM_ID_i_3_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_RAM_ID_i_4_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_RAM_ID_i_5_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_RAM_ID_i_6_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_RAM_ID_i_7_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_RAM_ID_i_8_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_RAM_ID_i_9_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_RAM_ID_i_10_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_RAM_ID_i_11_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_RAM_ID_i_12_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_RAM_ID_i_13_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_RAM_ID_i_14_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_RAM_ID_i_15_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_RAM_ID_i_16_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_RAM_ID_i_17_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_RAM_ID_i_18_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_RAM_ID_i_19_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_global_reset_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_scan_reset_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_RDATA_A1_o_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_RDATA_A1_o_1_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_RDATA_A1_o_2_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_RDATA_A1_o_3_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_RDATA_A1_o_4_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_RDATA_A1_o_5_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_RDATA_B1_o_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_RDATA_B1_o_1_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_RDATA_B1_o_2_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_RDATA_B1_o_3_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_RDATA_B1_o_4_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_RDATA_B1_o_5_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_RDATA_A1_o_6_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_RDATA_A1_o_7_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_RDATA_A1_o_8_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_RDATA_A1_o_9_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_RDATA_A1_o_10_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_RDATA_A1_o_11_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_RDATA_B1_o_6_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_RDATA_B1_o_7_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_RDATA_B1_o_8_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_RDATA_B1_o_9_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_RDATA_B1_o_10_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_1_subtile_0__pin_RDATA_B1_o_11_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_2_subtile_0__pin_RDATA_A1_o_12_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_2_subtile_0__pin_RDATA_A1_o_13_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_2_subtile_0__pin_RDATA_A1_o_14_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_2_subtile_0__pin_RDATA_A1_o_15_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_2_subtile_0__pin_RDATA_A1_o_16_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_2_subtile_0__pin_RDATA_A1_o_17_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_2_subtile_0__pin_RDATA_B1_o_12_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_2_subtile_0__pin_RDATA_B1_o_13_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_2_subtile_0__pin_RDATA_B1_o_14_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_2_subtile_0__pin_RDATA_B1_o_15_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_2_subtile_0__pin_RDATA_B1_o_16_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_2_subtile_0__pin_RDATA_B1_o_17_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_3_subtile_0__pin_RDATA_A2_o_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_3_subtile_0__pin_RDATA_A2_o_1_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_3_subtile_0__pin_RDATA_A2_o_2_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_3_subtile_0__pin_RDATA_A2_o_3_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_3_subtile_0__pin_RDATA_A2_o_4_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_3_subtile_0__pin_RDATA_A2_o_5_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_3_subtile_0__pin_RDATA_B2_o_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_3_subtile_0__pin_RDATA_B2_o_1_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_3_subtile_0__pin_RDATA_B2_o_2_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_3_subtile_0__pin_RDATA_B2_o_3_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_3_subtile_0__pin_RDATA_B2_o_4_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_3_subtile_0__pin_RDATA_B2_o_5_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_4_subtile_0__pin_RDATA_A2_o_6_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_4_subtile_0__pin_RDATA_A2_o_7_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_4_subtile_0__pin_RDATA_A2_o_8_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_4_subtile_0__pin_RDATA_A2_o_9_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_4_subtile_0__pin_RDATA_A2_o_10_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_4_subtile_0__pin_RDATA_A2_o_11_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_4_subtile_0__pin_RDATA_B2_o_6_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_4_subtile_0__pin_RDATA_B2_o_7_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_4_subtile_0__pin_RDATA_B2_o_8_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_4_subtile_0__pin_RDATA_B2_o_9_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_4_subtile_0__pin_RDATA_B2_o_10_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_4_subtile_0__pin_RDATA_B2_o_11_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_5_subtile_0__pin_RDATA_A2_o_12_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_5_subtile_0__pin_RDATA_A2_o_13_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_5_subtile_0__pin_RDATA_A2_o_14_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_5_subtile_0__pin_RDATA_A2_o_15_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_5_subtile_0__pin_RDATA_A2_o_16_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_5_subtile_0__pin_RDATA_A2_o_17_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_5_subtile_0__pin_RDATA_B2_o_12_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_5_subtile_0__pin_RDATA_B2_o_13_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_5_subtile_0__pin_RDATA_B2_o_14_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_5_subtile_0__pin_RDATA_B2_o_15_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_5_subtile_0__pin_RDATA_B2_o_16_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_5_subtile_0__pin_RDATA_B2_o_17_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_INIT_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ENA_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_REN_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_CLK_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_WEN_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_WEN_o_1_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_1_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_2_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_3_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_4_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_5_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_6_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_7_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_8_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_9_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_10_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_11_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_12_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_13_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_14_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_15_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_16_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_17_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_18_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_19_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_20_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_21_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_22_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_23_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_24_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_25_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_26_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_27_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_28_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_29_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_30_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_31_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_1_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_2_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_3_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_4_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_5_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_6_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_7_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_8_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_9_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_10_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_11_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_12_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_13_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_14_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_15_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_16_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_17_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_18_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_19_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_20_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_21_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_22_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_23_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_24_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_25_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_26_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_27_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_28_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_29_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_30_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_31_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_32_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_33_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_34_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_35_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_sc_out_1_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_sc_out_2_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_sc_out_3_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_sc_out_4_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_sc_out_5_;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	logical_tile_bram_mode_bram_ logical_tile_bram_mode_bram__0 (
		.test_en(test_en),
		.scan_mode(scan_mode),
		.scan_clk(scan_clk),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.bram_WDATA_A1_i({bottom_width_0_height_0_subtile_0__pin_WDATA_A1_i_0_, bottom_width_0_height_0_subtile_0__pin_WDATA_A1_i_1_, bottom_width_0_height_0_subtile_0__pin_WDATA_A1_i_2_, bottom_width_0_height_0_subtile_0__pin_WDATA_A1_i_3_, bottom_width_0_height_0_subtile_0__pin_WDATA_A1_i_4_, bottom_width_0_height_0_subtile_0__pin_WDATA_A1_i_5_, bottom_width_0_height_0_subtile_0__pin_WDATA_A1_i_6_, right_width_0_height_3_subtile_0__pin_WDATA_A1_i_7_, right_width_0_height_3_subtile_0__pin_WDATA_A1_i_8_, right_width_0_height_3_subtile_0__pin_WDATA_A1_i_9_, right_width_0_height_3_subtile_0__pin_WDATA_A1_i_10_, right_width_0_height_3_subtile_0__pin_WDATA_A1_i_11_, right_width_0_height_3_subtile_0__pin_WDATA_A1_i_12_, right_width_0_height_3_subtile_0__pin_WDATA_A1_i_13_, right_width_0_height_3_subtile_0__pin_WDATA_A1_i_14_, right_width_0_height_3_subtile_0__pin_WDATA_A1_i_15_, right_width_0_height_3_subtile_0__pin_WDATA_A1_i_16_, right_width_0_height_3_subtile_0__pin_WDATA_A1_i_17_}),
		.bram_WDATA_A2_i({right_width_0_height_4_subtile_0__pin_WDATA_A2_i_0_, right_width_0_height_4_subtile_0__pin_WDATA_A2_i_1_, right_width_0_height_4_subtile_0__pin_WDATA_A2_i_2_, right_width_0_height_4_subtile_0__pin_WDATA_A2_i_3_, right_width_0_height_4_subtile_0__pin_WDATA_A2_i_4_, right_width_0_height_4_subtile_0__pin_WDATA_A2_i_5_, right_width_0_height_4_subtile_0__pin_WDATA_A2_i_6_, right_width_0_height_4_subtile_0__pin_WDATA_A2_i_7_, right_width_0_height_4_subtile_0__pin_WDATA_A2_i_8_, right_width_0_height_2_subtile_0__pin_WDATA_A2_i_9_, right_width_0_height_2_subtile_0__pin_WDATA_A2_i_10_, right_width_0_height_2_subtile_0__pin_WDATA_A2_i_11_, right_width_0_height_2_subtile_0__pin_WDATA_A2_i_12_, right_width_0_height_2_subtile_0__pin_WDATA_A2_i_13_, right_width_0_height_2_subtile_0__pin_WDATA_A2_i_14_, right_width_0_height_2_subtile_0__pin_WDATA_A2_i_15_, right_width_0_height_2_subtile_0__pin_WDATA_A2_i_16_, right_width_0_height_1_subtile_0__pin_WDATA_A2_i_17_}),
		.bram_ADDR_A1_i({right_width_0_height_3_subtile_0__pin_ADDR_A1_i_0_, right_width_0_height_3_subtile_0__pin_ADDR_A1_i_1_, right_width_0_height_0_subtile_0__pin_ADDR_A1_i_2_, right_width_0_height_0_subtile_0__pin_ADDR_A1_i_3_, right_width_0_height_0_subtile_0__pin_ADDR_A1_i_4_, right_width_0_height_0_subtile_0__pin_ADDR_A1_i_5_, bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_6_, bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_7_, bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_8_, bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_9_, bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_10_, bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_11_, bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_12_, bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_13_, bottom_width_0_height_0_subtile_0__pin_ADDR_A1_i_14_}),
		.bram_ADDR_A2_i({right_width_0_height_2_subtile_0__pin_ADDR_A2_i_0_, right_width_0_height_1_subtile_0__pin_ADDR_A2_i_1_, right_width_0_height_2_subtile_0__pin_ADDR_A2_i_2_, right_width_0_height_2_subtile_0__pin_ADDR_A2_i_3_, right_width_0_height_2_subtile_0__pin_ADDR_A2_i_4_, right_width_0_height_2_subtile_0__pin_ADDR_A2_i_5_, right_width_0_height_2_subtile_0__pin_ADDR_A2_i_6_, right_width_0_height_2_subtile_0__pin_ADDR_A2_i_7_, right_width_0_height_2_subtile_0__pin_ADDR_A2_i_8_, right_width_0_height_2_subtile_0__pin_ADDR_A2_i_9_, right_width_0_height_2_subtile_0__pin_ADDR_A2_i_10_, right_width_0_height_2_subtile_0__pin_ADDR_A2_i_11_, right_width_0_height_2_subtile_0__pin_ADDR_A2_i_12_, right_width_0_height_2_subtile_0__pin_ADDR_A2_i_13_}),
		.bram_REN_A1_i(right_width_0_height_1_subtile_0__pin_REN_A1_i_0_),
		.bram_REN_A2_i(right_width_0_height_1_subtile_0__pin_REN_A2_i_0_),
		.bram_WEN_A1_i(right_width_0_height_2_subtile_0__pin_WEN_A1_i_0_),
		.bram_WEN_A2_i(right_width_0_height_1_subtile_0__pin_WEN_A2_i_0_),
		.bram_BE_A1_i({right_width_0_height_3_subtile_0__pin_BE_A1_i_0_, right_width_0_height_3_subtile_0__pin_BE_A1_i_1_}),
		.bram_BE_A2_i({right_width_0_height_1_subtile_0__pin_BE_A2_i_0_, right_width_0_height_1_subtile_0__pin_BE_A2_i_1_}),
		.bram_WDATA_B1_i({right_width_0_height_1_subtile_0__pin_WDATA_B1_i_0_, right_width_0_height_0_subtile_0__pin_WDATA_B1_i_1_, right_width_0_height_0_subtile_0__pin_WDATA_B1_i_2_, right_width_0_height_0_subtile_0__pin_WDATA_B1_i_3_, right_width_0_height_0_subtile_0__pin_WDATA_B1_i_4_, right_width_0_height_0_subtile_0__pin_WDATA_B1_i_5_, right_width_0_height_0_subtile_0__pin_WDATA_B1_i_6_, right_width_0_height_0_subtile_0__pin_WDATA_B1_i_7_, right_width_0_height_0_subtile_0__pin_WDATA_B1_i_8_, right_width_0_height_0_subtile_0__pin_WDATA_B1_i_9_, right_width_0_height_0_subtile_0__pin_WDATA_B1_i_10_, right_width_0_height_0_subtile_0__pin_WDATA_B1_i_11_, right_width_0_height_0_subtile_0__pin_WDATA_B1_i_12_, right_width_0_height_0_subtile_0__pin_WDATA_B1_i_13_, right_width_0_height_0_subtile_0__pin_WDATA_B1_i_14_, right_width_0_height_0_subtile_0__pin_WDATA_B1_i_15_, right_width_0_height_0_subtile_0__pin_WDATA_B1_i_16_, bottom_width_0_height_0_subtile_0__pin_WDATA_B1_i_17_}),
		.bram_WDATA_B2_i({right_width_0_height_5_subtile_0__pin_WDATA_B2_i_0_, right_width_0_height_5_subtile_0__pin_WDATA_B2_i_1_, right_width_0_height_5_subtile_0__pin_WDATA_B2_i_2_, right_width_0_height_5_subtile_0__pin_WDATA_B2_i_3_, right_width_0_height_5_subtile_0__pin_WDATA_B2_i_4_, right_width_0_height_5_subtile_0__pin_WDATA_B2_i_5_, right_width_0_height_5_subtile_0__pin_WDATA_B2_i_6_, right_width_0_height_5_subtile_0__pin_WDATA_B2_i_7_, right_width_0_height_5_subtile_0__pin_WDATA_B2_i_8_, right_width_0_height_5_subtile_0__pin_WDATA_B2_i_9_, right_width_0_height_5_subtile_0__pin_WDATA_B2_i_10_, right_width_0_height_5_subtile_0__pin_WDATA_B2_i_11_, right_width_0_height_5_subtile_0__pin_WDATA_B2_i_12_, right_width_0_height_5_subtile_0__pin_WDATA_B2_i_13_, right_width_0_height_5_subtile_0__pin_WDATA_B2_i_14_, right_width_0_height_5_subtile_0__pin_WDATA_B2_i_15_, right_width_0_height_5_subtile_0__pin_WDATA_B2_i_16_, right_width_0_height_4_subtile_0__pin_WDATA_B2_i_17_}),
		.bram_ADDR_B1_i({right_width_0_height_0_subtile_0__pin_ADDR_B1_i_0_, bottom_width_0_height_0_subtile_0__pin_ADDR_B1_i_1_, right_width_0_height_1_subtile_0__pin_ADDR_B1_i_2_, right_width_0_height_1_subtile_0__pin_ADDR_B1_i_3_, right_width_0_height_1_subtile_0__pin_ADDR_B1_i_4_, right_width_0_height_1_subtile_0__pin_ADDR_B1_i_5_, right_width_0_height_1_subtile_0__pin_ADDR_B1_i_6_, right_width_0_height_1_subtile_0__pin_ADDR_B1_i_7_, right_width_0_height_1_subtile_0__pin_ADDR_B1_i_8_, right_width_0_height_1_subtile_0__pin_ADDR_B1_i_9_, right_width_0_height_1_subtile_0__pin_ADDR_B1_i_10_, right_width_0_height_1_subtile_0__pin_ADDR_B1_i_11_, right_width_0_height_1_subtile_0__pin_ADDR_B1_i_12_, right_width_0_height_1_subtile_0__pin_ADDR_B1_i_13_, right_width_0_height_1_subtile_0__pin_ADDR_B1_i_14_}),
		.bram_ADDR_B2_i({right_width_0_height_5_subtile_0__pin_ADDR_B2_i_0_, right_width_0_height_4_subtile_0__pin_ADDR_B2_i_1_, right_width_0_height_5_subtile_0__pin_ADDR_B2_i_2_, right_width_0_height_5_subtile_0__pin_ADDR_B2_i_3_, right_width_0_height_4_subtile_0__pin_ADDR_B2_i_4_, right_width_0_height_4_subtile_0__pin_ADDR_B2_i_5_, right_width_0_height_4_subtile_0__pin_ADDR_B2_i_6_, right_width_0_height_4_subtile_0__pin_ADDR_B2_i_7_, right_width_0_height_4_subtile_0__pin_ADDR_B2_i_8_, right_width_0_height_4_subtile_0__pin_ADDR_B2_i_9_, right_width_0_height_4_subtile_0__pin_ADDR_B2_i_10_, right_width_0_height_4_subtile_0__pin_ADDR_B2_i_11_, right_width_0_height_4_subtile_0__pin_ADDR_B2_i_12_, right_width_0_height_4_subtile_0__pin_ADDR_B2_i_13_}),
		.bram_REN_B1_i(right_width_0_height_5_subtile_0__pin_REN_B1_i_0_),
		.bram_REN_B2_i(right_width_0_height_3_subtile_0__pin_REN_B2_i_0_),
		.bram_WEN_B1_i(right_width_0_height_4_subtile_0__pin_WEN_B1_i_0_),
		.bram_WEN_B2_i(right_width_0_height_3_subtile_0__pin_WEN_B2_i_0_),
		.bram_BE_B1_i({right_width_0_height_3_subtile_0__pin_BE_B1_i_0_, right_width_0_height_3_subtile_0__pin_BE_B1_i_1_}),
		.bram_BE_B2_i({right_width_0_height_3_subtile_0__pin_BE_B2_i_0_, right_width_0_height_3_subtile_0__pin_BE_B2_i_1_}),
		.bram_FLUSH1_i(right_width_0_height_3_subtile_0__pin_FLUSH1_i_0_),
		.bram_FLUSH2_i(right_width_0_height_1_subtile_0__pin_FLUSH2_i_0_),
		.bram_RAM_ID_i({left_width_0_height_0_subtile_0__pin_RAM_ID_i_0_, left_width_0_height_0_subtile_0__pin_RAM_ID_i_1_, left_width_0_height_0_subtile_0__pin_RAM_ID_i_2_, left_width_0_height_0_subtile_0__pin_RAM_ID_i_3_, left_width_0_height_0_subtile_0__pin_RAM_ID_i_4_, left_width_0_height_0_subtile_0__pin_RAM_ID_i_5_, left_width_0_height_0_subtile_0__pin_RAM_ID_i_6_, left_width_0_height_0_subtile_0__pin_RAM_ID_i_7_, left_width_0_height_0_subtile_0__pin_RAM_ID_i_8_, left_width_0_height_0_subtile_0__pin_RAM_ID_i_9_, left_width_0_height_0_subtile_0__pin_RAM_ID_i_10_, left_width_0_height_0_subtile_0__pin_RAM_ID_i_11_, left_width_0_height_0_subtile_0__pin_RAM_ID_i_12_, left_width_0_height_0_subtile_0__pin_RAM_ID_i_13_, left_width_0_height_0_subtile_0__pin_RAM_ID_i_14_, left_width_0_height_0_subtile_0__pin_RAM_ID_i_15_, left_width_0_height_0_subtile_0__pin_RAM_ID_i_16_, left_width_0_height_0_subtile_0__pin_RAM_ID_i_17_, left_width_0_height_0_subtile_0__pin_RAM_ID_i_18_, left_width_0_height_0_subtile_0__pin_RAM_ID_i_19_}),
		.bram_PL_INIT_i(top_width_0_height_0_subtile_0__pin_PL_INIT_i_0_),
		.bram_PL_ENA_i(top_width_0_height_0_subtile_0__pin_PL_ENA_i_0_),
		.bram_PL_REN_i(top_width_0_height_0_subtile_0__pin_PL_REN_i_0_),
		.bram_PL_WEN_i({top_width_0_height_0_subtile_0__pin_PL_WEN_i_0_, top_width_0_height_0_subtile_0__pin_PL_WEN_i_1_}),
		.bram_PL_ADDR_i({top_width_0_height_0_subtile_0__pin_PL_ADDR_i_0_, top_width_0_height_0_subtile_0__pin_PL_ADDR_i_1_, top_width_0_height_0_subtile_0__pin_PL_ADDR_i_2_, top_width_0_height_0_subtile_0__pin_PL_ADDR_i_3_, top_width_0_height_0_subtile_0__pin_PL_ADDR_i_4_, top_width_0_height_0_subtile_0__pin_PL_ADDR_i_5_, top_width_0_height_0_subtile_0__pin_PL_ADDR_i_6_, top_width_0_height_0_subtile_0__pin_PL_ADDR_i_7_, top_width_0_height_0_subtile_0__pin_PL_ADDR_i_8_, top_width_0_height_0_subtile_0__pin_PL_ADDR_i_9_, top_width_0_height_0_subtile_0__pin_PL_ADDR_i_10_, top_width_0_height_0_subtile_0__pin_PL_ADDR_i_11_, top_width_0_height_0_subtile_0__pin_PL_ADDR_i_12_, top_width_0_height_0_subtile_0__pin_PL_ADDR_i_13_, top_width_0_height_0_subtile_0__pin_PL_ADDR_i_14_, top_width_0_height_0_subtile_0__pin_PL_ADDR_i_15_, top_width_0_height_0_subtile_0__pin_PL_ADDR_i_16_, top_width_0_height_0_subtile_0__pin_PL_ADDR_i_17_, top_width_0_height_0_subtile_0__pin_PL_ADDR_i_18_, top_width_0_height_0_subtile_0__pin_PL_ADDR_i_19_, top_width_0_height_0_subtile_0__pin_PL_ADDR_i_20_, top_width_0_height_0_subtile_0__pin_PL_ADDR_i_21_, top_width_0_height_0_subtile_0__pin_PL_ADDR_i_22_, top_width_0_height_0_subtile_0__pin_PL_ADDR_i_23_, top_width_0_height_0_subtile_0__pin_PL_ADDR_i_24_, top_width_0_height_0_subtile_0__pin_PL_ADDR_i_25_, top_width_0_height_0_subtile_0__pin_PL_ADDR_i_26_, top_width_0_height_0_subtile_0__pin_PL_ADDR_i_27_, top_width_0_height_0_subtile_0__pin_PL_ADDR_i_28_, top_width_0_height_0_subtile_0__pin_PL_ADDR_i_29_, top_width_0_height_0_subtile_0__pin_PL_ADDR_i_30_, top_width_0_height_0_subtile_0__pin_PL_ADDR_i_31_}),
		.bram_PL_DATA_i({top_width_0_height_0_subtile_0__pin_PL_DATA_i_0_, top_width_0_height_0_subtile_0__pin_PL_DATA_i_1_, top_width_0_height_0_subtile_0__pin_PL_DATA_i_2_, top_width_0_height_0_subtile_0__pin_PL_DATA_i_3_, top_width_0_height_0_subtile_0__pin_PL_DATA_i_4_, top_width_0_height_0_subtile_0__pin_PL_DATA_i_5_, top_width_0_height_0_subtile_0__pin_PL_DATA_i_6_, top_width_0_height_0_subtile_0__pin_PL_DATA_i_7_, top_width_0_height_0_subtile_0__pin_PL_DATA_i_8_, top_width_0_height_0_subtile_0__pin_PL_DATA_i_9_, top_width_0_height_0_subtile_0__pin_PL_DATA_i_10_, top_width_0_height_0_subtile_0__pin_PL_DATA_i_11_, top_width_0_height_0_subtile_0__pin_PL_DATA_i_12_, top_width_0_height_0_subtile_0__pin_PL_DATA_i_13_, top_width_0_height_0_subtile_0__pin_PL_DATA_i_14_, top_width_0_height_0_subtile_0__pin_PL_DATA_i_15_, top_width_0_height_0_subtile_0__pin_PL_DATA_i_16_, top_width_0_height_0_subtile_0__pin_PL_DATA_i_17_, top_width_0_height_0_subtile_0__pin_PL_DATA_i_18_, top_width_0_height_0_subtile_0__pin_PL_DATA_i_19_, top_width_0_height_0_subtile_0__pin_PL_DATA_i_20_, top_width_0_height_0_subtile_0__pin_PL_DATA_i_21_, top_width_0_height_0_subtile_0__pin_PL_DATA_i_22_, top_width_0_height_0_subtile_0__pin_PL_DATA_i_23_, top_width_0_height_0_subtile_0__pin_PL_DATA_i_24_, top_width_0_height_0_subtile_0__pin_PL_DATA_i_25_, top_width_0_height_0_subtile_0__pin_PL_DATA_i_26_, top_width_0_height_0_subtile_0__pin_PL_DATA_i_27_, top_width_0_height_0_subtile_0__pin_PL_DATA_i_28_, top_width_0_height_0_subtile_0__pin_PL_DATA_i_29_, top_width_0_height_0_subtile_0__pin_PL_DATA_i_30_, top_width_0_height_0_subtile_0__pin_PL_DATA_i_31_, top_width_0_height_0_subtile_0__pin_PL_DATA_i_32_, top_width_0_height_0_subtile_0__pin_PL_DATA_i_33_, top_width_0_height_0_subtile_0__pin_PL_DATA_i_34_, top_width_0_height_0_subtile_0__pin_PL_DATA_i_35_}),
		.bram_global_reset(left_width_0_height_0_subtile_0__pin_global_reset_0_),
		.bram_scan_reset(left_width_0_height_0_subtile_0__pin_scan_reset_0_),
		.bram_sc_in({top_width_0_height_0_subtile_0__pin_sc_in_0_, top_width_0_height_0_subtile_0__pin_sc_in_1_, top_width_0_height_0_subtile_0__pin_sc_in_2_, top_width_0_height_0_subtile_0__pin_sc_in_3_, top_width_0_height_0_subtile_0__pin_sc_in_4_, top_width_0_height_0_subtile_0__pin_sc_in_5_}),
		.bram_PL_CLK_i(top_width_0_height_0_subtile_0__pin_PL_CLK_i_0_),
		.bram_clk({left_width_0_height_0_subtile_0__pin_clk_0_, left_width_0_height_0_subtile_0__pin_clk_1_, left_width_0_height_0_subtile_0__pin_clk_2_, left_width_0_height_0_subtile_0__pin_clk_3_}),
		.ccff_head(ccff_head),
		.bram_RDATA_A1_o({right_width_0_height_0_subtile_0__pin_RDATA_A1_o_0_, right_width_0_height_0_subtile_0__pin_RDATA_A1_o_1_, right_width_0_height_0_subtile_0__pin_RDATA_A1_o_2_, right_width_0_height_0_subtile_0__pin_RDATA_A1_o_3_, right_width_0_height_0_subtile_0__pin_RDATA_A1_o_4_, right_width_0_height_0_subtile_0__pin_RDATA_A1_o_5_, right_width_0_height_1_subtile_0__pin_RDATA_A1_o_6_, right_width_0_height_1_subtile_0__pin_RDATA_A1_o_7_, right_width_0_height_1_subtile_0__pin_RDATA_A1_o_8_, right_width_0_height_1_subtile_0__pin_RDATA_A1_o_9_, right_width_0_height_1_subtile_0__pin_RDATA_A1_o_10_, right_width_0_height_1_subtile_0__pin_RDATA_A1_o_11_, right_width_0_height_2_subtile_0__pin_RDATA_A1_o_12_, right_width_0_height_2_subtile_0__pin_RDATA_A1_o_13_, right_width_0_height_2_subtile_0__pin_RDATA_A1_o_14_, right_width_0_height_2_subtile_0__pin_RDATA_A1_o_15_, right_width_0_height_2_subtile_0__pin_RDATA_A1_o_16_, right_width_0_height_2_subtile_0__pin_RDATA_A1_o_17_}),
		.bram_RDATA_A2_o({right_width_0_height_3_subtile_0__pin_RDATA_A2_o_0_, right_width_0_height_3_subtile_0__pin_RDATA_A2_o_1_, right_width_0_height_3_subtile_0__pin_RDATA_A2_o_2_, right_width_0_height_3_subtile_0__pin_RDATA_A2_o_3_, right_width_0_height_3_subtile_0__pin_RDATA_A2_o_4_, right_width_0_height_3_subtile_0__pin_RDATA_A2_o_5_, right_width_0_height_4_subtile_0__pin_RDATA_A2_o_6_, right_width_0_height_4_subtile_0__pin_RDATA_A2_o_7_, right_width_0_height_4_subtile_0__pin_RDATA_A2_o_8_, right_width_0_height_4_subtile_0__pin_RDATA_A2_o_9_, right_width_0_height_4_subtile_0__pin_RDATA_A2_o_10_, right_width_0_height_4_subtile_0__pin_RDATA_A2_o_11_, right_width_0_height_5_subtile_0__pin_RDATA_A2_o_12_, right_width_0_height_5_subtile_0__pin_RDATA_A2_o_13_, right_width_0_height_5_subtile_0__pin_RDATA_A2_o_14_, right_width_0_height_5_subtile_0__pin_RDATA_A2_o_15_, right_width_0_height_5_subtile_0__pin_RDATA_A2_o_16_, right_width_0_height_5_subtile_0__pin_RDATA_A2_o_17_}),
		.bram_RDATA_B1_o({right_width_0_height_0_subtile_0__pin_RDATA_B1_o_0_, right_width_0_height_0_subtile_0__pin_RDATA_B1_o_1_, right_width_0_height_0_subtile_0__pin_RDATA_B1_o_2_, right_width_0_height_0_subtile_0__pin_RDATA_B1_o_3_, right_width_0_height_0_subtile_0__pin_RDATA_B1_o_4_, right_width_0_height_0_subtile_0__pin_RDATA_B1_o_5_, right_width_0_height_1_subtile_0__pin_RDATA_B1_o_6_, right_width_0_height_1_subtile_0__pin_RDATA_B1_o_7_, right_width_0_height_1_subtile_0__pin_RDATA_B1_o_8_, right_width_0_height_1_subtile_0__pin_RDATA_B1_o_9_, right_width_0_height_1_subtile_0__pin_RDATA_B1_o_10_, right_width_0_height_1_subtile_0__pin_RDATA_B1_o_11_, right_width_0_height_2_subtile_0__pin_RDATA_B1_o_12_, right_width_0_height_2_subtile_0__pin_RDATA_B1_o_13_, right_width_0_height_2_subtile_0__pin_RDATA_B1_o_14_, right_width_0_height_2_subtile_0__pin_RDATA_B1_o_15_, right_width_0_height_2_subtile_0__pin_RDATA_B1_o_16_, right_width_0_height_2_subtile_0__pin_RDATA_B1_o_17_}),
		.bram_RDATA_B2_o({right_width_0_height_3_subtile_0__pin_RDATA_B2_o_0_, right_width_0_height_3_subtile_0__pin_RDATA_B2_o_1_, right_width_0_height_3_subtile_0__pin_RDATA_B2_o_2_, right_width_0_height_3_subtile_0__pin_RDATA_B2_o_3_, right_width_0_height_3_subtile_0__pin_RDATA_B2_o_4_, right_width_0_height_3_subtile_0__pin_RDATA_B2_o_5_, right_width_0_height_4_subtile_0__pin_RDATA_B2_o_6_, right_width_0_height_4_subtile_0__pin_RDATA_B2_o_7_, right_width_0_height_4_subtile_0__pin_RDATA_B2_o_8_, right_width_0_height_4_subtile_0__pin_RDATA_B2_o_9_, right_width_0_height_4_subtile_0__pin_RDATA_B2_o_10_, right_width_0_height_4_subtile_0__pin_RDATA_B2_o_11_, right_width_0_height_5_subtile_0__pin_RDATA_B2_o_12_, right_width_0_height_5_subtile_0__pin_RDATA_B2_o_13_, right_width_0_height_5_subtile_0__pin_RDATA_B2_o_14_, right_width_0_height_5_subtile_0__pin_RDATA_B2_o_15_, right_width_0_height_5_subtile_0__pin_RDATA_B2_o_16_, right_width_0_height_5_subtile_0__pin_RDATA_B2_o_17_}),
		.bram_PL_INIT_o(bottom_width_0_height_0_subtile_0__pin_PL_INIT_o_0_),
		.bram_PL_ENA_o(bottom_width_0_height_0_subtile_0__pin_PL_ENA_o_0_),
		.bram_PL_REN_o(bottom_width_0_height_0_subtile_0__pin_PL_REN_o_0_),
		.bram_PL_CLK_o(bottom_width_0_height_0_subtile_0__pin_PL_CLK_o_0_),
		.bram_PL_WEN_o({bottom_width_0_height_0_subtile_0__pin_PL_WEN_o_0_, bottom_width_0_height_0_subtile_0__pin_PL_WEN_o_1_}),
		.bram_PL_ADDR_o({bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_0_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_1_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_2_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_3_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_4_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_5_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_6_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_7_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_8_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_9_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_10_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_11_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_12_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_13_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_14_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_15_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_16_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_17_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_18_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_19_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_20_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_21_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_22_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_23_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_24_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_25_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_26_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_27_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_28_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_29_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_30_, bottom_width_0_height_0_subtile_0__pin_PL_ADDR_o_31_}),
		.bram_PL_DATA_o({bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_0_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_1_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_2_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_3_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_4_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_5_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_6_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_7_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_8_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_9_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_10_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_11_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_12_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_13_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_14_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_15_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_16_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_17_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_18_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_19_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_20_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_21_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_22_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_23_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_24_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_25_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_26_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_27_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_28_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_29_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_30_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_31_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_32_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_33_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_34_, bottom_width_0_height_0_subtile_0__pin_PL_DATA_o_35_}),
		.bram_sc_out({bottom_width_0_height_0_subtile_0__pin_sc_out_0_, bottom_width_0_height_0_subtile_0__pin_sc_out_1_, bottom_width_0_height_0_subtile_0__pin_sc_out_2_, bottom_width_0_height_0_subtile_0__pin_sc_out_3_, bottom_width_0_height_0_subtile_0__pin_sc_out_4_, bottom_width_0_height_0_subtile_0__pin_sc_out_5_}),
		.ccff_tail(ccff_tail));

endmodule
// ----- END Verilog module for grid_bram -----

//----- Default net type -----
`default_nettype none



// ----- END Grid Verilog module: grid_bram -----

