// `timescale 1ns / 1ps

module and2(a,b,c);

input a, b;
output c;

assign c = a & b;

endmodule
