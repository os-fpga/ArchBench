//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for Unique Switch Blocks[0][8]
//	Author: Xifan TANG
//	Organization: University of Utah
//-------------------------------------------
//----- Time scale -----
`timescale 1ns / 1ps

//----- Default net type -----
`default_nettype wire

// ----- Verilog module for sb_0__8_ -----
module sb_0__8_(config_enable,
                prog_clock,
                chanx_right_in,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_8__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_9__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_10__pin_a2f_o_0_,
                right_bottom_grid_top_width_0_height_0_subtile_11__pin_a2f_o_0_,
                chany_bottom_in,
                bottom_right_grid_left_width_0_height_0_subtile_24__pin_a2f_o_0_,
                bottom_right_grid_left_width_0_height_0_subtile_25__pin_a2f_o_0_,
                bottom_right_grid_left_width_0_height_0_subtile_26__pin_a2f_o_0_,
                bottom_right_grid_left_width_0_height_0_subtile_27__pin_a2f_o_0_,
                bottom_right_grid_left_width_0_height_0_subtile_28__pin_a2f_o_0_,
                bottom_right_grid_left_width_0_height_0_subtile_29__pin_a2f_o_0_,
                bottom_right_grid_left_width_0_height_0_subtile_30__pin_a2f_o_0_,
                bottom_right_grid_left_width_0_height_0_subtile_31__pin_a2f_o_0_,
                bottom_right_grid_left_width_0_height_0_subtile_32__pin_a2f_o_0_,
                bottom_right_grid_left_width_0_height_0_subtile_33__pin_a2f_o_0_,
                bottom_right_grid_left_width_0_height_0_subtile_34__pin_a2f_o_0_,
                bottom_right_grid_left_width_0_height_0_subtile_35__pin_a2f_o_0_,
                bottom_right_grid_left_width_0_height_0_subtile_36__pin_a2f_o_0_,
                bottom_right_grid_left_width_0_height_0_subtile_37__pin_a2f_o_0_,
                bottom_right_grid_left_width_0_height_0_subtile_38__pin_a2f_o_0_,
                bottom_right_grid_left_width_0_height_0_subtile_39__pin_a2f_o_0_,
                bottom_right_grid_left_width_0_height_0_subtile_40__pin_a2f_o_0_,
                bottom_right_grid_left_width_0_height_0_subtile_41__pin_a2f_o_0_,
                bottom_right_grid_left_width_0_height_0_subtile_42__pin_a2f_o_0_,
                bottom_right_grid_left_width_0_height_0_subtile_43__pin_a2f_o_0_,
                bottom_right_grid_left_width_0_height_0_subtile_44__pin_a2f_o_0_,
                bottom_right_grid_left_width_0_height_0_subtile_45__pin_a2f_o_0_,
                bottom_right_grid_left_width_0_height_0_subtile_46__pin_a2f_o_0_,
                bottom_right_grid_left_width_0_height_0_subtile_47__pin_a2f_o_0_,
                bottom_right_grid_left_width_0_height_0_subtile_48__pin_a2f_o_0_,
                bottom_right_grid_left_width_0_height_0_subtile_49__pin_a2f_o_0_,
                bottom_right_grid_left_width_0_height_0_subtile_50__pin_a2f_o_0_,
                bottom_right_grid_left_width_0_height_0_subtile_51__pin_a2f_o_0_,
                bottom_right_grid_left_width_0_height_0_subtile_52__pin_a2f_o_0_,
                bottom_right_grid_left_width_0_height_0_subtile_53__pin_a2f_o_0_,
                bottom_right_grid_left_width_0_height_0_subtile_54__pin_a2f_o_0_,
                bottom_right_grid_left_width_0_height_0_subtile_55__pin_a2f_o_0_,
                bottom_right_grid_left_width_0_height_0_subtile_56__pin_a2f_o_0_,
                bottom_right_grid_left_width_0_height_0_subtile_57__pin_a2f_o_0_,
                bottom_right_grid_left_width_0_height_0_subtile_58__pin_a2f_o_0_,
                bottom_right_grid_left_width_0_height_0_subtile_59__pin_a2f_o_0_,
                bottom_right_grid_left_width_0_height_0_subtile_60__pin_a2f_o_0_,
                bottom_right_grid_left_width_0_height_0_subtile_61__pin_a2f_o_0_,
                bottom_right_grid_left_width_0_height_0_subtile_62__pin_a2f_o_0_,
                bottom_right_grid_left_width_0_height_0_subtile_63__pin_a2f_o_0_,
                bottom_right_grid_left_width_0_height_0_subtile_64__pin_a2f_o_0_,
                bottom_right_grid_left_width_0_height_0_subtile_65__pin_a2f_o_0_,
                bottom_right_grid_left_width_0_height_0_subtile_66__pin_a2f_o_0_,
                bottom_right_grid_left_width_0_height_0_subtile_67__pin_a2f_o_0_,
                bottom_right_grid_left_width_0_height_0_subtile_68__pin_a2f_o_0_,
                bottom_right_grid_left_width_0_height_0_subtile_69__pin_a2f_o_0_,
                bottom_right_grid_left_width_0_height_0_subtile_70__pin_a2f_o_0_,
                bottom_right_grid_left_width_0_height_0_subtile_71__pin_a2f_o_0_,
                ccff_head,
                chanx_right_out,
                chany_bottom_out,
                ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_clock;
//----- INPUT PORTS -----
input [0:95] chanx_right_in;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_8__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_9__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_10__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_11__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:95] chany_bottom_in;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_24__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_25__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_26__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_27__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_28__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_29__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_30__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_31__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_32__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_33__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_34__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_35__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_36__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_37__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_38__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_39__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_40__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_41__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_42__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_43__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_44__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_45__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_46__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_47__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_48__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_49__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_50__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_51__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_52__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_53__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_54__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_55__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_56__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_57__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_58__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_59__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_60__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_61__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_62__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_63__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_64__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_65__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_66__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_67__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_68__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_69__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_70__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_71__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:95] chanx_right_out;
//----- OUTPUT PORTS -----
output [0:95] chany_bottom_out;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:1] mux_tree_tapbuf_L2SB_size3_0_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size3_0_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size3_1_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size3_1_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size3_2_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size3_2_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size3_3_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size3_3_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size3_4_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size3_4_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size3_5_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size3_5_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size3_6_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size3_6_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size3_7_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size3_7_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size3_8_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size3_8_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_0_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_0_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_1_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_1_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_2_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_2_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_3_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_3_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_4_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_4_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_5_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_5_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_6_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_6_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_7_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_7_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_8_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_8_sram_inv;
wire [0:1] mux_tree_tapbuf_L2SB_size4_9_sram;
wire [0:1] mux_tree_tapbuf_L2SB_size4_9_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_0_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_0_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_10_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_10_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_11_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_11_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_12_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_12_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_13_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_13_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_14_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_14_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_15_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_15_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_16_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_16_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_17_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_17_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_18_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_18_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_19_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_19_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_1_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_1_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_20_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_20_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_21_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_21_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_22_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_22_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_23_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_23_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_24_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_24_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_25_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_25_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_26_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_26_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_27_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_27_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_28_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_28_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_29_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_29_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_2_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_2_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_30_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_30_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_31_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_31_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_32_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_32_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_33_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_33_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_34_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_34_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_35_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_35_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_36_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_36_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_37_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_37_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_38_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_38_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_39_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_39_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_3_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_3_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_40_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_40_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_41_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_41_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_42_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_42_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_43_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_43_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_44_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_44_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_45_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_45_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_46_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_46_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_47_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_47_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_48_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_48_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_49_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_49_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_4_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_4_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_50_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_50_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_51_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_51_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_52_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_52_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_53_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_53_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_54_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_54_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_5_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_5_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_6_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_6_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_7_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_7_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_8_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_8_sram_inv;
wire [0:1] mux_tree_tapbuf_L4SB_size3_9_sram;
wire [0:1] mux_tree_tapbuf_L4SB_size3_9_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_0_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_0_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_10_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_10_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_1_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_1_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_2_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_2_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_3_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_3_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_4_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_4_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_5_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_5_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_6_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_6_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_7_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_7_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_8_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_8_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size7_9_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size7_9_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_0_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_0_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_10_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_10_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_11_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_11_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_12_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_12_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_13_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_13_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_14_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_14_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_15_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_15_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_16_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_16_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_17_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_17_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_18_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_18_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_19_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_19_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_1_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_1_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_20_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_20_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_21_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_21_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_22_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_22_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_23_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_23_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_24_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_24_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_25_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_25_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_26_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_26_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_27_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_27_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_28_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_28_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_29_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_29_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_2_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_2_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_30_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_30_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_31_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_31_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_32_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_32_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_33_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_33_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_34_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_34_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_35_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_35_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_36_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_36_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_37_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_37_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_38_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_38_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_39_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_39_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_3_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_3_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_40_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_40_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_41_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_41_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_42_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_42_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_43_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_43_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_44_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_44_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_45_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_45_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_46_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_46_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_47_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_47_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_48_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_48_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_49_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_49_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_4_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_4_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_50_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_50_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_51_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_51_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_52_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_52_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_53_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_53_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_54_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_54_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_55_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_55_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_56_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_56_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_57_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_57_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_58_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_58_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_59_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_59_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_5_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_5_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_60_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_60_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_61_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_61_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_62_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_62_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_63_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_63_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_64_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_64_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_65_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_65_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_6_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_6_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_7_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_7_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_8_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_8_sram_inv;
wire [0:2] mux_tree_tapbuf_L4SB_size8_9_sram;
wire [0:2] mux_tree_tapbuf_L4SB_size8_9_sram_inv;

// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 184 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[18] = chany_bottom_in[76];
// ----- Local connection due to Wire 185 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[17] = chany_bottom_in[77];
// ----- Local connection due to Wire 186 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[16] = chany_bottom_in[78];
// ----- Local connection due to Wire 187 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[15] = chany_bottom_in[79];
// ----- Local connection due to Wire 188 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[14] = chany_bottom_in[80];
// ----- Local connection due to Wire 189 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[13] = chany_bottom_in[81];
// ----- Local connection due to Wire 190 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[12] = chany_bottom_in[82];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	mux_tree_tapbuf_L2SB_size2 mux_right_track_0 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, chany_bottom_in[94]}),
		.sram(mux_tree_tapbuf_L2SB_size2_0_sram),
		.sram_inv(mux_tree_tapbuf_L2SB_size2_0_sram_inv),
		.out(chanx_right_out[0]));

	mux_tree_tapbuf_L2SB_size2 mux_right_track_2 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, chany_bottom_in[93]}),
		.sram(mux_tree_tapbuf_L2SB_size2_1_sram),
		.sram_inv(mux_tree_tapbuf_L2SB_size2_1_sram_inv),
		.out(chanx_right_out[1]));

	mux_tree_tapbuf_L2SB_size2 mux_right_track_4 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, chany_bottom_in[92]}),
		.sram(mux_tree_tapbuf_L2SB_size2_2_sram),
		.sram_inv(mux_tree_tapbuf_L2SB_size2_2_sram_inv),
		.out(chanx_right_out[2]));

	mux_tree_tapbuf_L2SB_size2 mux_right_track_6 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, chany_bottom_in[91]}),
		.sram(mux_tree_tapbuf_L2SB_size2_3_sram),
		.sram_inv(mux_tree_tapbuf_L2SB_size2_3_sram_inv),
		.out(chanx_right_out[3]));

	mux_tree_tapbuf_L2SB_size2 mux_right_track_8 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_, chany_bottom_in[90]}),
		.sram(mux_tree_tapbuf_L2SB_size2_4_sram),
		.sram_inv(mux_tree_tapbuf_L2SB_size2_4_sram_inv),
		.out(chanx_right_out[4]));

	mux_tree_tapbuf_L2SB_size2 mux_right_track_10 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_, chany_bottom_in[89]}),
		.sram(mux_tree_tapbuf_L2SB_size2_5_sram),
		.sram_inv(mux_tree_tapbuf_L2SB_size2_5_sram_inv),
		.out(chanx_right_out[5]));

	mux_tree_tapbuf_L2SB_size2 mux_right_track_12 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_, chany_bottom_in[88]}),
		.sram(mux_tree_tapbuf_L2SB_size2_6_sram),
		.sram_inv(mux_tree_tapbuf_L2SB_size2_6_sram_inv),
		.out(chanx_right_out[6]));

	mux_tree_tapbuf_L2SB_size2 mux_right_track_14 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_, chany_bottom_in[87]}),
		.sram(mux_tree_tapbuf_L2SB_size2_7_sram),
		.sram_inv(mux_tree_tapbuf_L2SB_size2_7_sram_inv),
		.out(chanx_right_out[7]));

	mux_tree_tapbuf_L2SB_size2 mux_right_track_16 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_8__pin_a2f_o_0_, chany_bottom_in[86]}),
		.sram(mux_tree_tapbuf_L2SB_size2_8_sram),
		.sram_inv(mux_tree_tapbuf_L2SB_size2_8_sram_inv),
		.out(chanx_right_out[8]));

	mux_tree_tapbuf_L2SB_size2 mux_right_track_18 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_9__pin_a2f_o_0_, chany_bottom_in[85]}),
		.sram(mux_tree_tapbuf_L2SB_size2_9_sram),
		.sram_inv(mux_tree_tapbuf_L2SB_size2_9_sram_inv),
		.out(chanx_right_out[9]));

	mux_tree_tapbuf_L2SB_size2 mux_right_track_20 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_10__pin_a2f_o_0_, chany_bottom_in[84]}),
		.sram(mux_tree_tapbuf_L2SB_size2_10_sram),
		.sram_inv(mux_tree_tapbuf_L2SB_size2_10_sram_inv),
		.out(chanx_right_out[10]));

	mux_tree_tapbuf_L2SB_size2 mux_right_track_22 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_11__pin_a2f_o_0_, chany_bottom_in[83]}),
		.sram(mux_tree_tapbuf_L2SB_size2_11_sram),
		.sram_inv(mux_tree_tapbuf_L2SB_size2_11_sram_inv),
		.out(chanx_right_out[11]));

	mux_tree_tapbuf_L2SB_size2_mem mem_right_track_0 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(ccff_head),
		.ccff_tail(mux_tree_tapbuf_L2SB_size2_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size2_0_sram),
		.mem_outb(mux_tree_tapbuf_L2SB_size2_0_sram_inv));

	mux_tree_tapbuf_L2SB_size2_mem mem_right_track_2 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size2_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size2_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size2_1_sram),
		.mem_outb(mux_tree_tapbuf_L2SB_size2_1_sram_inv));

	mux_tree_tapbuf_L2SB_size2_mem mem_right_track_4 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size2_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size2_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size2_2_sram),
		.mem_outb(mux_tree_tapbuf_L2SB_size2_2_sram_inv));

	mux_tree_tapbuf_L2SB_size2_mem mem_right_track_6 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size2_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size2_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size2_3_sram),
		.mem_outb(mux_tree_tapbuf_L2SB_size2_3_sram_inv));

	mux_tree_tapbuf_L2SB_size2_mem mem_right_track_8 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size2_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size2_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size2_4_sram),
		.mem_outb(mux_tree_tapbuf_L2SB_size2_4_sram_inv));

	mux_tree_tapbuf_L2SB_size2_mem mem_right_track_10 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size2_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size2_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size2_5_sram),
		.mem_outb(mux_tree_tapbuf_L2SB_size2_5_sram_inv));

	mux_tree_tapbuf_L2SB_size2_mem mem_right_track_12 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size2_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size2_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size2_6_sram),
		.mem_outb(mux_tree_tapbuf_L2SB_size2_6_sram_inv));

	mux_tree_tapbuf_L2SB_size2_mem mem_right_track_14 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size2_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size2_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size2_7_sram),
		.mem_outb(mux_tree_tapbuf_L2SB_size2_7_sram_inv));

	mux_tree_tapbuf_L2SB_size2_mem mem_right_track_16 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size2_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size2_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size2_8_sram),
		.mem_outb(mux_tree_tapbuf_L2SB_size2_8_sram_inv));

	mux_tree_tapbuf_L2SB_size2_mem mem_right_track_18 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size2_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size2_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size2_9_sram),
		.mem_outb(mux_tree_tapbuf_L2SB_size2_9_sram_inv));

	mux_tree_tapbuf_L2SB_size2_mem mem_right_track_20 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size2_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size2_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size2_10_sram),
		.mem_outb(mux_tree_tapbuf_L2SB_size2_10_sram_inv));

	mux_tree_tapbuf_L2SB_size2_mem mem_right_track_22 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size2_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size2_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size2_11_sram),
		.mem_outb(mux_tree_tapbuf_L2SB_size2_11_sram_inv));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_38 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_, chany_bottom_in[75]}),
		.sram(mux_tree_tapbuf_L4SB_size3_0_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_0_sram_inv[0:1]),
		.out(chanx_right_out[19]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_40 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_8__pin_a2f_o_0_, chany_bottom_in[74]}),
		.sram(mux_tree_tapbuf_L4SB_size3_1_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_1_sram_inv[0:1]),
		.out(chanx_right_out[20]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_42 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_9__pin_a2f_o_0_, chany_bottom_in[73]}),
		.sram(mux_tree_tapbuf_L4SB_size3_2_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_2_sram_inv[0:1]),
		.out(chanx_right_out[21]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_44 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_10__pin_a2f_o_0_, chany_bottom_in[72]}),
		.sram(mux_tree_tapbuf_L4SB_size3_3_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_3_sram_inv[0:1]),
		.out(chanx_right_out[22]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_46 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_11__pin_a2f_o_0_, chany_bottom_in[71]}),
		.sram(mux_tree_tapbuf_L4SB_size3_4_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_4_sram_inv[0:1]),
		.out(chanx_right_out[23]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_52 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_, chany_bottom_in[68]}),
		.sram(mux_tree_tapbuf_L4SB_size3_5_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_5_sram_inv[0:1]),
		.out(chanx_right_out[26]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_54 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_8__pin_a2f_o_0_, chany_bottom_in[67]}),
		.sram(mux_tree_tapbuf_L4SB_size3_6_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_6_sram_inv[0:1]),
		.out(chanx_right_out[27]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_56 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_9__pin_a2f_o_0_, chany_bottom_in[66]}),
		.sram(mux_tree_tapbuf_L4SB_size3_7_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_7_sram_inv[0:1]),
		.out(chanx_right_out[28]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_58 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_10__pin_a2f_o_0_, chany_bottom_in[65]}),
		.sram(mux_tree_tapbuf_L4SB_size3_8_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_8_sram_inv[0:1]),
		.out(chanx_right_out[29]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_60 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_11__pin_a2f_o_0_, chany_bottom_in[64]}),
		.sram(mux_tree_tapbuf_L4SB_size3_9_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_9_sram_inv[0:1]),
		.out(chanx_right_out[30]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_66 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_, chany_bottom_in[61]}),
		.sram(mux_tree_tapbuf_L4SB_size3_10_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_10_sram_inv[0:1]),
		.out(chanx_right_out[33]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_68 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_8__pin_a2f_o_0_, chany_bottom_in[60]}),
		.sram(mux_tree_tapbuf_L4SB_size3_11_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_11_sram_inv[0:1]),
		.out(chanx_right_out[34]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_70 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_9__pin_a2f_o_0_, chany_bottom_in[59]}),
		.sram(mux_tree_tapbuf_L4SB_size3_12_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_12_sram_inv[0:1]),
		.out(chanx_right_out[35]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_72 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_10__pin_a2f_o_0_, chany_bottom_in[58]}),
		.sram(mux_tree_tapbuf_L4SB_size3_13_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_13_sram_inv[0:1]),
		.out(chanx_right_out[36]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_74 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_11__pin_a2f_o_0_, chany_bottom_in[57]}),
		.sram(mux_tree_tapbuf_L4SB_size3_14_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_14_sram_inv[0:1]),
		.out(chanx_right_out[37]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_80 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_, chany_bottom_in[54]}),
		.sram(mux_tree_tapbuf_L4SB_size3_15_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_15_sram_inv[0:1]),
		.out(chanx_right_out[40]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_82 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_8__pin_a2f_o_0_, chany_bottom_in[53]}),
		.sram(mux_tree_tapbuf_L4SB_size3_16_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_16_sram_inv[0:1]),
		.out(chanx_right_out[41]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_84 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_9__pin_a2f_o_0_, chany_bottom_in[52]}),
		.sram(mux_tree_tapbuf_L4SB_size3_17_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_17_sram_inv[0:1]),
		.out(chanx_right_out[42]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_86 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_10__pin_a2f_o_0_, chany_bottom_in[51]}),
		.sram(mux_tree_tapbuf_L4SB_size3_18_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_18_sram_inv[0:1]),
		.out(chanx_right_out[43]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_88 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_11__pin_a2f_o_0_, chany_bottom_in[50]}),
		.sram(mux_tree_tapbuf_L4SB_size3_19_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_19_sram_inv[0:1]),
		.out(chanx_right_out[44]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_94 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_, chany_bottom_in[47]}),
		.sram(mux_tree_tapbuf_L4SB_size3_20_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_20_sram_inv[0:1]),
		.out(chanx_right_out[47]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_96 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_8__pin_a2f_o_0_, chany_bottom_in[46]}),
		.sram(mux_tree_tapbuf_L4SB_size3_21_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_21_sram_inv[0:1]),
		.out(chanx_right_out[48]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_98 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_9__pin_a2f_o_0_, chany_bottom_in[45]}),
		.sram(mux_tree_tapbuf_L4SB_size3_22_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_22_sram_inv[0:1]),
		.out(chanx_right_out[49]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_100 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_10__pin_a2f_o_0_, chany_bottom_in[44]}),
		.sram(mux_tree_tapbuf_L4SB_size3_23_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_23_sram_inv[0:1]),
		.out(chanx_right_out[50]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_102 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_11__pin_a2f_o_0_, chany_bottom_in[43]}),
		.sram(mux_tree_tapbuf_L4SB_size3_24_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_24_sram_inv[0:1]),
		.out(chanx_right_out[51]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_108 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_, chany_bottom_in[40]}),
		.sram(mux_tree_tapbuf_L4SB_size3_25_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_25_sram_inv[0:1]),
		.out(chanx_right_out[54]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_110 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_8__pin_a2f_o_0_, chany_bottom_in[39]}),
		.sram(mux_tree_tapbuf_L4SB_size3_26_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_26_sram_inv[0:1]),
		.out(chanx_right_out[55]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_112 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_9__pin_a2f_o_0_, chany_bottom_in[38]}),
		.sram(mux_tree_tapbuf_L4SB_size3_27_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_27_sram_inv[0:1]),
		.out(chanx_right_out[56]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_114 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_10__pin_a2f_o_0_, chany_bottom_in[37]}),
		.sram(mux_tree_tapbuf_L4SB_size3_28_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_28_sram_inv[0:1]),
		.out(chanx_right_out[57]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_116 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_11__pin_a2f_o_0_, chany_bottom_in[36]}),
		.sram(mux_tree_tapbuf_L4SB_size3_29_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_29_sram_inv[0:1]),
		.out(chanx_right_out[58]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_122 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_, chany_bottom_in[33]}),
		.sram(mux_tree_tapbuf_L4SB_size3_30_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_30_sram_inv[0:1]),
		.out(chanx_right_out[61]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_124 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_8__pin_a2f_o_0_, chany_bottom_in[32]}),
		.sram(mux_tree_tapbuf_L4SB_size3_31_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_31_sram_inv[0:1]),
		.out(chanx_right_out[62]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_126 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_9__pin_a2f_o_0_, chany_bottom_in[31]}),
		.sram(mux_tree_tapbuf_L4SB_size3_32_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_32_sram_inv[0:1]),
		.out(chanx_right_out[63]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_128 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_10__pin_a2f_o_0_, chany_bottom_in[30]}),
		.sram(mux_tree_tapbuf_L4SB_size3_33_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_33_sram_inv[0:1]),
		.out(chanx_right_out[64]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_130 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_11__pin_a2f_o_0_, chany_bottom_in[29]}),
		.sram(mux_tree_tapbuf_L4SB_size3_34_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_34_sram_inv[0:1]),
		.out(chanx_right_out[65]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_136 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_, chany_bottom_in[26]}),
		.sram(mux_tree_tapbuf_L4SB_size3_35_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_35_sram_inv[0:1]),
		.out(chanx_right_out[68]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_138 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_8__pin_a2f_o_0_, chany_bottom_in[25]}),
		.sram(mux_tree_tapbuf_L4SB_size3_36_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_36_sram_inv[0:1]),
		.out(chanx_right_out[69]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_140 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_9__pin_a2f_o_0_, chany_bottom_in[24]}),
		.sram(mux_tree_tapbuf_L4SB_size3_37_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_37_sram_inv[0:1]),
		.out(chanx_right_out[70]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_142 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_10__pin_a2f_o_0_, chany_bottom_in[23]}),
		.sram(mux_tree_tapbuf_L4SB_size3_38_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_38_sram_inv[0:1]),
		.out(chanx_right_out[71]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_144 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_11__pin_a2f_o_0_, chany_bottom_in[22]}),
		.sram(mux_tree_tapbuf_L4SB_size3_39_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_39_sram_inv[0:1]),
		.out(chanx_right_out[72]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_150 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_, chany_bottom_in[19]}),
		.sram(mux_tree_tapbuf_L4SB_size3_40_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_40_sram_inv[0:1]),
		.out(chanx_right_out[75]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_152 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_8__pin_a2f_o_0_, chany_bottom_in[18]}),
		.sram(mux_tree_tapbuf_L4SB_size3_41_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_41_sram_inv[0:1]),
		.out(chanx_right_out[76]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_154 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_9__pin_a2f_o_0_, chany_bottom_in[17]}),
		.sram(mux_tree_tapbuf_L4SB_size3_42_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_42_sram_inv[0:1]),
		.out(chanx_right_out[77]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_156 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_10__pin_a2f_o_0_, chany_bottom_in[16]}),
		.sram(mux_tree_tapbuf_L4SB_size3_43_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_43_sram_inv[0:1]),
		.out(chanx_right_out[78]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_158 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_11__pin_a2f_o_0_, chany_bottom_in[15]}),
		.sram(mux_tree_tapbuf_L4SB_size3_44_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_44_sram_inv[0:1]),
		.out(chanx_right_out[79]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_164 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_, chany_bottom_in[12]}),
		.sram(mux_tree_tapbuf_L4SB_size3_45_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_45_sram_inv[0:1]),
		.out(chanx_right_out[82]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_166 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_8__pin_a2f_o_0_, chany_bottom_in[11]}),
		.sram(mux_tree_tapbuf_L4SB_size3_46_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_46_sram_inv[0:1]),
		.out(chanx_right_out[83]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_168 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_9__pin_a2f_o_0_, chany_bottom_in[10]}),
		.sram(mux_tree_tapbuf_L4SB_size3_47_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_47_sram_inv[0:1]),
		.out(chanx_right_out[84]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_170 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_10__pin_a2f_o_0_, chany_bottom_in[9]}),
		.sram(mux_tree_tapbuf_L4SB_size3_48_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_48_sram_inv[0:1]),
		.out(chanx_right_out[85]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_172 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_11__pin_a2f_o_0_, chany_bottom_in[8]}),
		.sram(mux_tree_tapbuf_L4SB_size3_49_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_49_sram_inv[0:1]),
		.out(chanx_right_out[86]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_178 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_, chany_bottom_in[5]}),
		.sram(mux_tree_tapbuf_L4SB_size3_50_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_50_sram_inv[0:1]),
		.out(chanx_right_out[89]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_180 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_8__pin_a2f_o_0_, chany_bottom_in[4]}),
		.sram(mux_tree_tapbuf_L4SB_size3_51_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_51_sram_inv[0:1]),
		.out(chanx_right_out[90]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_182 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_9__pin_a2f_o_0_, chany_bottom_in[3]}),
		.sram(mux_tree_tapbuf_L4SB_size3_52_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_52_sram_inv[0:1]),
		.out(chanx_right_out[91]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_184 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_10__pin_a2f_o_0_, chany_bottom_in[2]}),
		.sram(mux_tree_tapbuf_L4SB_size3_53_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_53_sram_inv[0:1]),
		.out(chanx_right_out[92]));

	mux_tree_tapbuf_L4SB_size3 mux_right_track_186 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_11__pin_a2f_o_0_, chany_bottom_in[1]}),
		.sram(mux_tree_tapbuf_L4SB_size3_54_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L4SB_size3_54_sram_inv[0:1]),
		.out(chanx_right_out[93]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_38 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size2_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_0_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_0_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_40 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_1_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_1_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_42 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_2_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_2_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_44 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_3_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_3_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_46 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_4_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_4_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_52 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size2_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_5_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_5_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_54 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_6_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_6_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_56 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_7_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_7_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_58 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_8_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_8_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_60 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_9_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_9_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_66 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size2_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_10_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_10_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_68 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_11_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_11_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_70 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_12_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_12_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_72 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_13_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_13_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_74 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_14_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_14_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_80 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size2_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_15_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_15_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_82 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_16_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_16_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_84 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_17_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_17_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_86 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_18_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_18_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_88 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_19_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_19_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_94 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size2_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_20_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_20_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_96 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_21_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_21_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_98 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_22_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_22_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_100 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_23_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_23_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_102 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_24_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_24_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_108 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size2_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_25_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_25_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_110 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_26_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_26_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_112 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_27_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_27_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_27_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_114 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_27_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_28_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_28_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_28_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_116 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_28_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_29_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_29_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_29_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_122 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size2_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_30_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_30_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_30_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_124 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_30_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_31_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_31_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_31_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_126 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_31_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_32_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_32_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_32_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_128 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_32_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_33_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_33_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_33_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_130 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_33_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_34_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_34_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_34_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_136 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size2_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_35_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_35_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_35_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_138 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_35_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_36_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_36_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_36_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_140 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_36_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_37_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_37_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_37_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_142 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_37_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_38_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_38_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_38_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_144 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_38_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_39_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_39_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_39_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_150 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size2_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_40_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_40_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_40_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_152 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_40_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_41_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_41_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_41_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_154 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_41_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_42_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_42_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_42_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_156 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_42_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_43_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_43_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_43_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_158 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_43_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_44_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_44_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_44_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_164 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size2_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_45_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_45_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_45_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_166 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_45_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_46_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_46_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_46_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_168 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_46_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_47_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_47_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_47_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_170 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_47_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_48_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_48_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_48_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_172 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_48_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_49_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_49_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_49_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_178 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size2_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_50_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_50_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_50_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_180 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_50_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_51_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_51_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_51_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_182 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_51_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_52_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_52_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_52_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_184 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_52_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_53_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_53_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_53_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size3_mem mem_right_track_186 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_53_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size3_mem_54_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size3_54_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L4SB_size3_54_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size2 mux_right_track_48 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_, chany_bottom_in[70]}),
		.sram(mux_tree_tapbuf_L4SB_size2_0_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_0_sram_inv),
		.out(chanx_right_out[24]));

	mux_tree_tapbuf_L4SB_size2 mux_right_track_50 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_, chany_bottom_in[69]}),
		.sram(mux_tree_tapbuf_L4SB_size2_1_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_1_sram_inv),
		.out(chanx_right_out[25]));

	mux_tree_tapbuf_L4SB_size2 mux_right_track_62 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_, chany_bottom_in[63]}),
		.sram(mux_tree_tapbuf_L4SB_size2_2_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_2_sram_inv),
		.out(chanx_right_out[31]));

	mux_tree_tapbuf_L4SB_size2 mux_right_track_64 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_, chany_bottom_in[62]}),
		.sram(mux_tree_tapbuf_L4SB_size2_3_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_3_sram_inv),
		.out(chanx_right_out[32]));

	mux_tree_tapbuf_L4SB_size2 mux_right_track_76 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_, chany_bottom_in[56]}),
		.sram(mux_tree_tapbuf_L4SB_size2_4_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_4_sram_inv),
		.out(chanx_right_out[38]));

	mux_tree_tapbuf_L4SB_size2 mux_right_track_78 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_, chany_bottom_in[55]}),
		.sram(mux_tree_tapbuf_L4SB_size2_5_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_5_sram_inv),
		.out(chanx_right_out[39]));

	mux_tree_tapbuf_L4SB_size2 mux_right_track_90 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_, chany_bottom_in[49]}),
		.sram(mux_tree_tapbuf_L4SB_size2_6_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_6_sram_inv),
		.out(chanx_right_out[45]));

	mux_tree_tapbuf_L4SB_size2 mux_right_track_92 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_, chany_bottom_in[48]}),
		.sram(mux_tree_tapbuf_L4SB_size2_7_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_7_sram_inv),
		.out(chanx_right_out[46]));

	mux_tree_tapbuf_L4SB_size2 mux_right_track_104 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_, chany_bottom_in[42]}),
		.sram(mux_tree_tapbuf_L4SB_size2_8_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_8_sram_inv),
		.out(chanx_right_out[52]));

	mux_tree_tapbuf_L4SB_size2 mux_right_track_106 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_, chany_bottom_in[41]}),
		.sram(mux_tree_tapbuf_L4SB_size2_9_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_9_sram_inv),
		.out(chanx_right_out[53]));

	mux_tree_tapbuf_L4SB_size2 mux_right_track_118 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_, chany_bottom_in[35]}),
		.sram(mux_tree_tapbuf_L4SB_size2_10_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_10_sram_inv),
		.out(chanx_right_out[59]));

	mux_tree_tapbuf_L4SB_size2 mux_right_track_120 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_, chany_bottom_in[34]}),
		.sram(mux_tree_tapbuf_L4SB_size2_11_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_11_sram_inv),
		.out(chanx_right_out[60]));

	mux_tree_tapbuf_L4SB_size2 mux_right_track_132 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_, chany_bottom_in[28]}),
		.sram(mux_tree_tapbuf_L4SB_size2_12_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_12_sram_inv),
		.out(chanx_right_out[66]));

	mux_tree_tapbuf_L4SB_size2 mux_right_track_134 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_, chany_bottom_in[27]}),
		.sram(mux_tree_tapbuf_L4SB_size2_13_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_13_sram_inv),
		.out(chanx_right_out[67]));

	mux_tree_tapbuf_L4SB_size2 mux_right_track_146 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_, chany_bottom_in[21]}),
		.sram(mux_tree_tapbuf_L4SB_size2_14_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_14_sram_inv),
		.out(chanx_right_out[73]));

	mux_tree_tapbuf_L4SB_size2 mux_right_track_148 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_, chany_bottom_in[20]}),
		.sram(mux_tree_tapbuf_L4SB_size2_15_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_15_sram_inv),
		.out(chanx_right_out[74]));

	mux_tree_tapbuf_L4SB_size2 mux_right_track_160 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_, chany_bottom_in[14]}),
		.sram(mux_tree_tapbuf_L4SB_size2_16_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_16_sram_inv),
		.out(chanx_right_out[80]));

	mux_tree_tapbuf_L4SB_size2 mux_right_track_162 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_, chany_bottom_in[13]}),
		.sram(mux_tree_tapbuf_L4SB_size2_17_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_17_sram_inv),
		.out(chanx_right_out[81]));

	mux_tree_tapbuf_L4SB_size2 mux_right_track_174 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_, chany_bottom_in[7]}),
		.sram(mux_tree_tapbuf_L4SB_size2_18_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_18_sram_inv),
		.out(chanx_right_out[87]));

	mux_tree_tapbuf_L4SB_size2 mux_right_track_176 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_, chany_bottom_in[6]}),
		.sram(mux_tree_tapbuf_L4SB_size2_19_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_19_sram_inv),
		.out(chanx_right_out[88]));

	mux_tree_tapbuf_L4SB_size2 mux_right_track_188 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_, chany_bottom_in[0]}),
		.sram(mux_tree_tapbuf_L4SB_size2_20_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_20_sram_inv),
		.out(chanx_right_out[94]));

	mux_tree_tapbuf_L4SB_size2 mux_right_track_190 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_, chany_bottom_in[95]}),
		.sram(mux_tree_tapbuf_L4SB_size2_21_sram),
		.sram_inv(mux_tree_tapbuf_L4SB_size2_21_sram_inv),
		.out(chanx_right_out[95]));

	mux_tree_tapbuf_L4SB_size2_mem mem_right_track_48 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size2_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size2_0_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_0_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_right_track_50 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size2_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size2_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size2_1_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_1_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_right_track_62 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size2_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size2_2_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_2_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_right_track_64 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size2_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size2_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size2_3_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_3_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_right_track_76 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size2_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size2_4_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_4_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_right_track_78 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size2_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size2_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size2_5_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_5_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_right_track_90 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size2_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size2_6_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_6_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_right_track_92 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size2_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size2_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size2_7_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_7_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_right_track_104 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size2_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size2_8_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_8_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_right_track_106 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size2_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size2_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size2_9_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_9_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_right_track_118 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_29_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size2_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size2_10_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_10_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_right_track_120 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size2_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size2_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size2_11_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_11_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_right_track_132 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_34_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size2_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size2_12_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_12_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_right_track_134 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size2_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size2_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size2_13_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_13_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_right_track_146 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_39_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size2_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size2_14_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_14_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_right_track_148 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size2_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size2_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size2_15_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_15_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_right_track_160 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_44_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size2_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size2_16_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_16_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_right_track_162 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size2_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size2_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size2_17_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_17_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_right_track_174 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_49_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size2_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size2_18_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_18_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_right_track_176 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size2_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size2_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size2_19_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_19_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_right_track_188 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size3_mem_54_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size2_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size2_20_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_20_sram_inv));

	mux_tree_tapbuf_L4SB_size2_mem mem_right_track_190 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size2_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size2_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size2_21_sram),
		.mem_outb(mux_tree_tapbuf_L4SB_size2_21_sram_inv));

	mux_tree_tapbuf_L2SB_size4 mux_bottom_track_1 (
		.in({chanx_right_in[94], bottom_right_grid_left_width_0_height_0_subtile_24__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_43__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_62__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L2SB_size4_0_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_0_sram_inv[0:1]),
		.out(chany_bottom_out[0]));

	mux_tree_tapbuf_L2SB_size4 mux_bottom_track_3 (
		.in({chanx_right_in[93], bottom_right_grid_left_width_0_height_0_subtile_25__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_44__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_63__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L2SB_size4_1_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_1_sram_inv[0:1]),
		.out(chany_bottom_out[1]));

	mux_tree_tapbuf_L2SB_size4 mux_bottom_track_5 (
		.in({chanx_right_in[92], bottom_right_grid_left_width_0_height_0_subtile_26__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_45__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_64__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L2SB_size4_2_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_2_sram_inv[0:1]),
		.out(chany_bottom_out[2]));

	mux_tree_tapbuf_L2SB_size4 mux_bottom_track_7 (
		.in({chanx_right_in[91], bottom_right_grid_left_width_0_height_0_subtile_27__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_46__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_65__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L2SB_size4_3_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_3_sram_inv[0:1]),
		.out(chany_bottom_out[3]));

	mux_tree_tapbuf_L2SB_size4 mux_bottom_track_9 (
		.in({chanx_right_in[90], bottom_right_grid_left_width_0_height_0_subtile_28__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_47__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_66__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L2SB_size4_4_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_4_sram_inv[0:1]),
		.out(chany_bottom_out[4]));

	mux_tree_tapbuf_L2SB_size4 mux_bottom_track_11 (
		.in({chanx_right_in[89], bottom_right_grid_left_width_0_height_0_subtile_29__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_48__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_67__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L2SB_size4_5_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_5_sram_inv[0:1]),
		.out(chany_bottom_out[5]));

	mux_tree_tapbuf_L2SB_size4 mux_bottom_track_13 (
		.in({chanx_right_in[88], bottom_right_grid_left_width_0_height_0_subtile_30__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_49__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_68__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L2SB_size4_6_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_6_sram_inv[0:1]),
		.out(chany_bottom_out[6]));

	mux_tree_tapbuf_L2SB_size4 mux_bottom_track_15 (
		.in({chanx_right_in[87], bottom_right_grid_left_width_0_height_0_subtile_31__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_50__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_69__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L2SB_size4_7_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_7_sram_inv[0:1]),
		.out(chany_bottom_out[7]));

	mux_tree_tapbuf_L2SB_size4 mux_bottom_track_17 (
		.in({chanx_right_in[86], bottom_right_grid_left_width_0_height_0_subtile_32__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_51__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_70__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L2SB_size4_8_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_8_sram_inv[0:1]),
		.out(chany_bottom_out[8]));

	mux_tree_tapbuf_L2SB_size4 mux_bottom_track_19 (
		.in({chanx_right_in[85], bottom_right_grid_left_width_0_height_0_subtile_33__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_52__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_71__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L2SB_size4_9_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size4_9_sram_inv[0:1]),
		.out(chany_bottom_out[9]));

	mux_tree_tapbuf_L2SB_size4_mem mem_bottom_track_1 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size2_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_0_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_0_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_bottom_track_3 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_1_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_1_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_bottom_track_5 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_2_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_2_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_bottom_track_7 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_3_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_3_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_bottom_track_9 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_4_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_4_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_bottom_track_11 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_5_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_5_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_bottom_track_13 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_6_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_6_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_bottom_track_15 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_7_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_7_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_bottom_track_17 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_8_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_8_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size4_mem mem_bottom_track_19 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size4_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size4_9_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size4_9_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size3 mux_bottom_track_21 (
		.in({chanx_right_in[84], bottom_right_grid_left_width_0_height_0_subtile_34__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_53__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L2SB_size3_0_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size3_0_sram_inv[0:1]),
		.out(chany_bottom_out[10]));

	mux_tree_tapbuf_L2SB_size3 mux_bottom_track_23 (
		.in({chanx_right_in[83], bottom_right_grid_left_width_0_height_0_subtile_35__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_54__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L2SB_size3_1_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size3_1_sram_inv[0:1]),
		.out(chany_bottom_out[11]));

	mux_tree_tapbuf_L2SB_size3 mux_bottom_track_25 (
		.in({chanx_right_in[82], bottom_right_grid_left_width_0_height_0_subtile_36__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_55__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L2SB_size3_2_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size3_2_sram_inv[0:1]),
		.out(chany_bottom_out[12]));

	mux_tree_tapbuf_L2SB_size3 mux_bottom_track_27 (
		.in({chanx_right_in[81], bottom_right_grid_left_width_0_height_0_subtile_37__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_56__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L2SB_size3_3_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size3_3_sram_inv[0:1]),
		.out(chany_bottom_out[13]));

	mux_tree_tapbuf_L2SB_size3 mux_bottom_track_29 (
		.in({chanx_right_in[80], bottom_right_grid_left_width_0_height_0_subtile_38__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_57__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L2SB_size3_4_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size3_4_sram_inv[0:1]),
		.out(chany_bottom_out[14]));

	mux_tree_tapbuf_L2SB_size3 mux_bottom_track_31 (
		.in({chanx_right_in[79], bottom_right_grid_left_width_0_height_0_subtile_39__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_58__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L2SB_size3_5_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size3_5_sram_inv[0:1]),
		.out(chany_bottom_out[15]));

	mux_tree_tapbuf_L2SB_size3 mux_bottom_track_33 (
		.in({chanx_right_in[78], bottom_right_grid_left_width_0_height_0_subtile_40__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_59__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L2SB_size3_6_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size3_6_sram_inv[0:1]),
		.out(chany_bottom_out[16]));

	mux_tree_tapbuf_L2SB_size3 mux_bottom_track_35 (
		.in({chanx_right_in[77], bottom_right_grid_left_width_0_height_0_subtile_41__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_60__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L2SB_size3_7_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size3_7_sram_inv[0:1]),
		.out(chany_bottom_out[17]));

	mux_tree_tapbuf_L2SB_size3 mux_bottom_track_37 (
		.in({chanx_right_in[76], bottom_right_grid_left_width_0_height_0_subtile_42__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_61__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L2SB_size3_8_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_L2SB_size3_8_sram_inv[0:1]),
		.out(chany_bottom_out[18]));

	mux_tree_tapbuf_L2SB_size3_mem mem_bottom_track_21 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size4_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size3_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size3_0_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size3_0_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size3_mem mem_bottom_track_23 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size3_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size3_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size3_1_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size3_1_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size3_mem mem_bottom_track_25 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size3_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size3_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size3_2_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size3_2_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size3_mem mem_bottom_track_27 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size3_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size3_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size3_3_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size3_3_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size3_mem mem_bottom_track_29 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size3_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size3_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size3_4_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size3_4_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size3_mem mem_bottom_track_31 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size3_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size3_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size3_5_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size3_5_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size3_mem mem_bottom_track_33 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size3_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size3_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size3_6_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size3_6_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size3_mem mem_bottom_track_35 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size3_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size3_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size3_7_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size3_7_sram_inv[0:1]));

	mux_tree_tapbuf_L2SB_size3_mem mem_bottom_track_37 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size3_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L2SB_size3_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_L2SB_size3_8_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_L2SB_size3_8_sram_inv[0:1]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_39 (
		.in({chanx_right_in[75], bottom_right_grid_left_width_0_height_0_subtile_24__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_31__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_38__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_45__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_52__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_59__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_66__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_0_sram_inv[0:2]),
		.out(chany_bottom_out[19]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_41 (
		.in({chanx_right_in[74], bottom_right_grid_left_width_0_height_0_subtile_25__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_32__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_39__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_46__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_53__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_60__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_67__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_1_sram_inv[0:2]),
		.out(chany_bottom_out[20]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_43 (
		.in({chanx_right_in[73], bottom_right_grid_left_width_0_height_0_subtile_26__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_33__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_40__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_47__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_54__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_61__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_68__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_2_sram_inv[0:2]),
		.out(chany_bottom_out[21]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_45 (
		.in({chanx_right_in[72], bottom_right_grid_left_width_0_height_0_subtile_27__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_34__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_41__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_48__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_55__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_62__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_69__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_3_sram_inv[0:2]),
		.out(chany_bottom_out[22]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_47 (
		.in({chanx_right_in[71], bottom_right_grid_left_width_0_height_0_subtile_28__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_35__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_42__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_49__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_56__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_63__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_70__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_4_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_4_sram_inv[0:2]),
		.out(chany_bottom_out[23]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_49 (
		.in({chanx_right_in[70], bottom_right_grid_left_width_0_height_0_subtile_29__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_36__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_43__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_50__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_57__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_64__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_71__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_5_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_5_sram_inv[0:2]),
		.out(chany_bottom_out[24]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_53 (
		.in({chanx_right_in[68], bottom_right_grid_left_width_0_height_0_subtile_24__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_31__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_38__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_45__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_52__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_59__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_66__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_6_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_6_sram_inv[0:2]),
		.out(chany_bottom_out[26]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_55 (
		.in({chanx_right_in[67], bottom_right_grid_left_width_0_height_0_subtile_25__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_32__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_39__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_46__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_53__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_60__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_67__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_7_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_7_sram_inv[0:2]),
		.out(chany_bottom_out[27]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_57 (
		.in({chanx_right_in[66], bottom_right_grid_left_width_0_height_0_subtile_26__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_33__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_40__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_47__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_54__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_61__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_68__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_8_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_8_sram_inv[0:2]),
		.out(chany_bottom_out[28]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_59 (
		.in({chanx_right_in[65], bottom_right_grid_left_width_0_height_0_subtile_27__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_34__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_41__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_48__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_55__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_62__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_69__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_9_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_9_sram_inv[0:2]),
		.out(chany_bottom_out[29]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_61 (
		.in({chanx_right_in[64], bottom_right_grid_left_width_0_height_0_subtile_28__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_35__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_42__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_49__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_56__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_63__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_70__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_10_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_10_sram_inv[0:2]),
		.out(chany_bottom_out[30]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_63 (
		.in({chanx_right_in[63], bottom_right_grid_left_width_0_height_0_subtile_29__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_36__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_43__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_50__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_57__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_64__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_71__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_11_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_11_sram_inv[0:2]),
		.out(chany_bottom_out[31]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_67 (
		.in({chanx_right_in[61], bottom_right_grid_left_width_0_height_0_subtile_24__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_31__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_38__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_45__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_52__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_59__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_66__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_12_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_12_sram_inv[0:2]),
		.out(chany_bottom_out[33]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_69 (
		.in({chanx_right_in[60], bottom_right_grid_left_width_0_height_0_subtile_25__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_32__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_39__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_46__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_53__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_60__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_67__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_13_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_13_sram_inv[0:2]),
		.out(chany_bottom_out[34]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_71 (
		.in({chanx_right_in[59], bottom_right_grid_left_width_0_height_0_subtile_26__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_33__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_40__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_47__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_54__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_61__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_68__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_14_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_14_sram_inv[0:2]),
		.out(chany_bottom_out[35]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_73 (
		.in({chanx_right_in[58], bottom_right_grid_left_width_0_height_0_subtile_27__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_34__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_41__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_48__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_55__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_62__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_69__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_15_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_15_sram_inv[0:2]),
		.out(chany_bottom_out[36]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_75 (
		.in({chanx_right_in[57], bottom_right_grid_left_width_0_height_0_subtile_28__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_35__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_42__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_49__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_56__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_63__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_70__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_16_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_16_sram_inv[0:2]),
		.out(chany_bottom_out[37]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_77 (
		.in({chanx_right_in[56], bottom_right_grid_left_width_0_height_0_subtile_29__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_36__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_43__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_50__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_57__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_64__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_71__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_17_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_17_sram_inv[0:2]),
		.out(chany_bottom_out[38]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_81 (
		.in({chanx_right_in[54], bottom_right_grid_left_width_0_height_0_subtile_24__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_31__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_38__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_45__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_52__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_59__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_66__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_18_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_18_sram_inv[0:2]),
		.out(chany_bottom_out[40]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_83 (
		.in({chanx_right_in[53], bottom_right_grid_left_width_0_height_0_subtile_25__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_32__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_39__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_46__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_53__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_60__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_67__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_19_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_19_sram_inv[0:2]),
		.out(chany_bottom_out[41]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_85 (
		.in({chanx_right_in[52], bottom_right_grid_left_width_0_height_0_subtile_26__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_33__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_40__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_47__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_54__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_61__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_68__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_20_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_20_sram_inv[0:2]),
		.out(chany_bottom_out[42]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_87 (
		.in({chanx_right_in[51], bottom_right_grid_left_width_0_height_0_subtile_27__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_34__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_41__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_48__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_55__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_62__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_69__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_21_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_21_sram_inv[0:2]),
		.out(chany_bottom_out[43]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_89 (
		.in({chanx_right_in[50], bottom_right_grid_left_width_0_height_0_subtile_28__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_35__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_42__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_49__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_56__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_63__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_70__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_22_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_22_sram_inv[0:2]),
		.out(chany_bottom_out[44]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_91 (
		.in({chanx_right_in[49], bottom_right_grid_left_width_0_height_0_subtile_29__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_36__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_43__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_50__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_57__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_64__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_71__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_23_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_23_sram_inv[0:2]),
		.out(chany_bottom_out[45]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_95 (
		.in({chanx_right_in[47], bottom_right_grid_left_width_0_height_0_subtile_24__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_31__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_38__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_45__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_52__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_59__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_66__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_24_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_24_sram_inv[0:2]),
		.out(chany_bottom_out[47]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_97 (
		.in({chanx_right_in[46], bottom_right_grid_left_width_0_height_0_subtile_25__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_32__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_39__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_46__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_53__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_60__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_67__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_25_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_25_sram_inv[0:2]),
		.out(chany_bottom_out[48]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_99 (
		.in({chanx_right_in[45], bottom_right_grid_left_width_0_height_0_subtile_26__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_33__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_40__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_47__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_54__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_61__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_68__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_26_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_26_sram_inv[0:2]),
		.out(chany_bottom_out[49]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_101 (
		.in({chanx_right_in[44], bottom_right_grid_left_width_0_height_0_subtile_27__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_34__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_41__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_48__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_55__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_62__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_69__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_27_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_27_sram_inv[0:2]),
		.out(chany_bottom_out[50]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_103 (
		.in({chanx_right_in[43], bottom_right_grid_left_width_0_height_0_subtile_28__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_35__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_42__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_49__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_56__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_63__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_70__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_28_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_28_sram_inv[0:2]),
		.out(chany_bottom_out[51]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_105 (
		.in({chanx_right_in[42], bottom_right_grid_left_width_0_height_0_subtile_29__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_36__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_43__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_50__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_57__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_64__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_71__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_29_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_29_sram_inv[0:2]),
		.out(chany_bottom_out[52]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_109 (
		.in({chanx_right_in[40], bottom_right_grid_left_width_0_height_0_subtile_24__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_31__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_38__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_45__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_52__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_59__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_66__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_30_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_30_sram_inv[0:2]),
		.out(chany_bottom_out[54]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_111 (
		.in({chanx_right_in[39], bottom_right_grid_left_width_0_height_0_subtile_25__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_32__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_39__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_46__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_53__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_60__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_67__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_31_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_31_sram_inv[0:2]),
		.out(chany_bottom_out[55]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_113 (
		.in({chanx_right_in[38], bottom_right_grid_left_width_0_height_0_subtile_26__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_33__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_40__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_47__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_54__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_61__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_68__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_32_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_32_sram_inv[0:2]),
		.out(chany_bottom_out[56]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_115 (
		.in({chanx_right_in[37], bottom_right_grid_left_width_0_height_0_subtile_27__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_34__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_41__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_48__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_55__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_62__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_69__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_33_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_33_sram_inv[0:2]),
		.out(chany_bottom_out[57]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_117 (
		.in({chanx_right_in[36], bottom_right_grid_left_width_0_height_0_subtile_28__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_35__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_42__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_49__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_56__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_63__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_70__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_34_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_34_sram_inv[0:2]),
		.out(chany_bottom_out[58]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_119 (
		.in({chanx_right_in[35], bottom_right_grid_left_width_0_height_0_subtile_29__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_36__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_43__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_50__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_57__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_64__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_71__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_35_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_35_sram_inv[0:2]),
		.out(chany_bottom_out[59]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_123 (
		.in({chanx_right_in[33], bottom_right_grid_left_width_0_height_0_subtile_24__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_31__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_38__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_45__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_52__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_59__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_66__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_36_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_36_sram_inv[0:2]),
		.out(chany_bottom_out[61]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_125 (
		.in({chanx_right_in[32], bottom_right_grid_left_width_0_height_0_subtile_25__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_32__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_39__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_46__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_53__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_60__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_67__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_37_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_37_sram_inv[0:2]),
		.out(chany_bottom_out[62]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_127 (
		.in({chanx_right_in[31], bottom_right_grid_left_width_0_height_0_subtile_26__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_33__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_40__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_47__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_54__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_61__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_68__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_38_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_38_sram_inv[0:2]),
		.out(chany_bottom_out[63]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_129 (
		.in({chanx_right_in[30], bottom_right_grid_left_width_0_height_0_subtile_27__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_34__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_41__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_48__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_55__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_62__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_69__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_39_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_39_sram_inv[0:2]),
		.out(chany_bottom_out[64]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_131 (
		.in({chanx_right_in[29], bottom_right_grid_left_width_0_height_0_subtile_28__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_35__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_42__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_49__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_56__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_63__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_70__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_40_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_40_sram_inv[0:2]),
		.out(chany_bottom_out[65]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_133 (
		.in({chanx_right_in[28], bottom_right_grid_left_width_0_height_0_subtile_29__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_36__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_43__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_50__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_57__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_64__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_71__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_41_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_41_sram_inv[0:2]),
		.out(chany_bottom_out[66]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_137 (
		.in({chanx_right_in[26], bottom_right_grid_left_width_0_height_0_subtile_24__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_31__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_38__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_45__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_52__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_59__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_66__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_42_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_42_sram_inv[0:2]),
		.out(chany_bottom_out[68]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_139 (
		.in({chanx_right_in[25], bottom_right_grid_left_width_0_height_0_subtile_25__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_32__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_39__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_46__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_53__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_60__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_67__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_43_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_43_sram_inv[0:2]),
		.out(chany_bottom_out[69]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_141 (
		.in({chanx_right_in[24], bottom_right_grid_left_width_0_height_0_subtile_26__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_33__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_40__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_47__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_54__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_61__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_68__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_44_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_44_sram_inv[0:2]),
		.out(chany_bottom_out[70]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_143 (
		.in({chanx_right_in[23], bottom_right_grid_left_width_0_height_0_subtile_27__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_34__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_41__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_48__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_55__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_62__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_69__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_45_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_45_sram_inv[0:2]),
		.out(chany_bottom_out[71]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_145 (
		.in({chanx_right_in[22], bottom_right_grid_left_width_0_height_0_subtile_28__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_35__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_42__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_49__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_56__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_63__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_70__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_46_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_46_sram_inv[0:2]),
		.out(chany_bottom_out[72]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_147 (
		.in({chanx_right_in[21], bottom_right_grid_left_width_0_height_0_subtile_29__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_36__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_43__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_50__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_57__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_64__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_71__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_47_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_47_sram_inv[0:2]),
		.out(chany_bottom_out[73]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_151 (
		.in({chanx_right_in[19], bottom_right_grid_left_width_0_height_0_subtile_24__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_31__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_38__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_45__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_52__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_59__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_66__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_48_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_48_sram_inv[0:2]),
		.out(chany_bottom_out[75]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_153 (
		.in({chanx_right_in[18], bottom_right_grid_left_width_0_height_0_subtile_25__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_32__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_39__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_46__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_53__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_60__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_67__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_49_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_49_sram_inv[0:2]),
		.out(chany_bottom_out[76]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_155 (
		.in({chanx_right_in[17], bottom_right_grid_left_width_0_height_0_subtile_26__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_33__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_40__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_47__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_54__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_61__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_68__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_50_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_50_sram_inv[0:2]),
		.out(chany_bottom_out[77]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_157 (
		.in({chanx_right_in[16], bottom_right_grid_left_width_0_height_0_subtile_27__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_34__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_41__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_48__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_55__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_62__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_69__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_51_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_51_sram_inv[0:2]),
		.out(chany_bottom_out[78]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_159 (
		.in({chanx_right_in[15], bottom_right_grid_left_width_0_height_0_subtile_28__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_35__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_42__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_49__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_56__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_63__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_70__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_52_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_52_sram_inv[0:2]),
		.out(chany_bottom_out[79]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_161 (
		.in({chanx_right_in[14], bottom_right_grid_left_width_0_height_0_subtile_29__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_36__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_43__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_50__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_57__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_64__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_71__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_53_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_53_sram_inv[0:2]),
		.out(chany_bottom_out[80]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_165 (
		.in({chanx_right_in[12], bottom_right_grid_left_width_0_height_0_subtile_24__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_31__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_38__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_45__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_52__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_59__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_66__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_54_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_54_sram_inv[0:2]),
		.out(chany_bottom_out[82]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_167 (
		.in({chanx_right_in[11], bottom_right_grid_left_width_0_height_0_subtile_25__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_32__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_39__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_46__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_53__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_60__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_67__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_55_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_55_sram_inv[0:2]),
		.out(chany_bottom_out[83]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_169 (
		.in({chanx_right_in[10], bottom_right_grid_left_width_0_height_0_subtile_26__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_33__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_40__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_47__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_54__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_61__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_68__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_56_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_56_sram_inv[0:2]),
		.out(chany_bottom_out[84]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_171 (
		.in({chanx_right_in[9], bottom_right_grid_left_width_0_height_0_subtile_27__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_34__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_41__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_48__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_55__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_62__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_69__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_57_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_57_sram_inv[0:2]),
		.out(chany_bottom_out[85]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_173 (
		.in({chanx_right_in[8], bottom_right_grid_left_width_0_height_0_subtile_28__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_35__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_42__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_49__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_56__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_63__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_70__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_58_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_58_sram_inv[0:2]),
		.out(chany_bottom_out[86]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_175 (
		.in({chanx_right_in[7], bottom_right_grid_left_width_0_height_0_subtile_29__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_36__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_43__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_50__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_57__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_64__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_71__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_59_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_59_sram_inv[0:2]),
		.out(chany_bottom_out[87]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_179 (
		.in({chanx_right_in[5], bottom_right_grid_left_width_0_height_0_subtile_24__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_31__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_38__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_45__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_52__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_59__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_66__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_60_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_60_sram_inv[0:2]),
		.out(chany_bottom_out[89]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_181 (
		.in({chanx_right_in[4], bottom_right_grid_left_width_0_height_0_subtile_25__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_32__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_39__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_46__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_53__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_60__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_67__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_61_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_61_sram_inv[0:2]),
		.out(chany_bottom_out[90]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_183 (
		.in({chanx_right_in[3], bottom_right_grid_left_width_0_height_0_subtile_26__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_33__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_40__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_47__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_54__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_61__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_68__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_62_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_62_sram_inv[0:2]),
		.out(chany_bottom_out[91]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_185 (
		.in({chanx_right_in[2], bottom_right_grid_left_width_0_height_0_subtile_27__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_34__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_41__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_48__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_55__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_62__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_69__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_63_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_63_sram_inv[0:2]),
		.out(chany_bottom_out[92]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_187 (
		.in({chanx_right_in[1], bottom_right_grid_left_width_0_height_0_subtile_28__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_35__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_42__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_49__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_56__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_63__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_70__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_64_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_64_sram_inv[0:2]),
		.out(chany_bottom_out[93]));

	mux_tree_tapbuf_L4SB_size8 mux_bottom_track_189 (
		.in({chanx_right_in[0], bottom_right_grid_left_width_0_height_0_subtile_29__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_36__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_43__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_50__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_57__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_64__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_71__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size8_65_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size8_65_sram_inv[0:2]),
		.out(chany_bottom_out[94]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_39 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L2SB_size3_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_0_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_41 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_1_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_43 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_2_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_45 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_3_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_47 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_4_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_4_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_49 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_5_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_5_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_53 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size7_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_6_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_6_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_55 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_7_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_7_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_57 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_8_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_8_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_59 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_9_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_9_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_61 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_10_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_10_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_63 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_11_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_11_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_67 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size7_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_12_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_12_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_69 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_13_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_13_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_71 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_14_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_14_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_73 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_15_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_15_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_75 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_16_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_16_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_77 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_17_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_17_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_81 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size7_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_18_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_18_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_83 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_19_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_19_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_85 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_20_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_20_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_87 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_21_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_21_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_89 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_22_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_22_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_91 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_23_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_23_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_95 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size7_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_24_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_24_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_97 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_25_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_25_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_99 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_26_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_26_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_101 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_27_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_27_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_27_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_103 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_27_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_28_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_28_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_28_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_105 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_28_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_29_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_29_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_29_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_109 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size7_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_30_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_30_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_30_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_111 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_30_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_31_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_31_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_31_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_113 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_31_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_32_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_32_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_32_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_115 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_32_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_33_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_33_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_33_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_117 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_33_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_34_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_34_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_34_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_119 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_34_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_35_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_35_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_35_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_123 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size7_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_36_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_36_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_36_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_125 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_36_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_37_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_37_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_37_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_127 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_37_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_38_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_38_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_38_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_129 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_38_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_39_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_39_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_39_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_131 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_39_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_40_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_40_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_40_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_133 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_40_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_41_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_41_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_41_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_137 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size7_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_42_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_42_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_42_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_139 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_42_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_43_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_43_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_43_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_141 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_43_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_44_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_44_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_44_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_143 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_44_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_45_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_45_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_45_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_145 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_45_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_46_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_46_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_46_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_147 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_46_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_47_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_47_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_47_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_151 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size7_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_48_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_48_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_48_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_153 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_48_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_49_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_49_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_49_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_155 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_49_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_50_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_50_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_50_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_157 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_50_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_51_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_51_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_51_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_159 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_51_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_52_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_52_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_52_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_161 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_52_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_53_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_53_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_53_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_165 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size7_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_54_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_54_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_54_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_167 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_54_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_55_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_55_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_55_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_169 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_55_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_56_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_56_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_56_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_171 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_56_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_57_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_57_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_57_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_173 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_57_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_58_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_58_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_58_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_175 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_58_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_59_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_59_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_59_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_179 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size7_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_60_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_60_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_60_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_181 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_60_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_61_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_61_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_61_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_183 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_61_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_62_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_62_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_62_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_185 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_62_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_63_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_63_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_63_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_187 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_63_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_64_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_64_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_64_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size8_mem mem_bottom_track_189 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_64_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size8_mem_65_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size8_65_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size8_65_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7 mux_bottom_track_51 (
		.in({chanx_right_in[69], bottom_right_grid_left_width_0_height_0_subtile_30__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_37__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_44__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_51__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_58__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_65__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size7_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_0_sram_inv[0:2]),
		.out(chany_bottom_out[25]));

	mux_tree_tapbuf_L4SB_size7 mux_bottom_track_65 (
		.in({chanx_right_in[62], bottom_right_grid_left_width_0_height_0_subtile_30__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_37__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_44__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_51__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_58__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_65__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size7_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_1_sram_inv[0:2]),
		.out(chany_bottom_out[32]));

	mux_tree_tapbuf_L4SB_size7 mux_bottom_track_79 (
		.in({chanx_right_in[55], bottom_right_grid_left_width_0_height_0_subtile_30__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_37__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_44__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_51__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_58__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_65__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size7_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_2_sram_inv[0:2]),
		.out(chany_bottom_out[39]));

	mux_tree_tapbuf_L4SB_size7 mux_bottom_track_93 (
		.in({chanx_right_in[48], bottom_right_grid_left_width_0_height_0_subtile_30__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_37__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_44__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_51__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_58__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_65__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size7_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_3_sram_inv[0:2]),
		.out(chany_bottom_out[46]));

	mux_tree_tapbuf_L4SB_size7 mux_bottom_track_107 (
		.in({chanx_right_in[41], bottom_right_grid_left_width_0_height_0_subtile_30__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_37__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_44__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_51__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_58__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_65__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size7_4_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_4_sram_inv[0:2]),
		.out(chany_bottom_out[53]));

	mux_tree_tapbuf_L4SB_size7 mux_bottom_track_121 (
		.in({chanx_right_in[34], bottom_right_grid_left_width_0_height_0_subtile_30__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_37__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_44__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_51__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_58__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_65__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size7_5_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_5_sram_inv[0:2]),
		.out(chany_bottom_out[60]));

	mux_tree_tapbuf_L4SB_size7 mux_bottom_track_135 (
		.in({chanx_right_in[27], bottom_right_grid_left_width_0_height_0_subtile_30__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_37__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_44__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_51__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_58__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_65__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size7_6_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_6_sram_inv[0:2]),
		.out(chany_bottom_out[67]));

	mux_tree_tapbuf_L4SB_size7 mux_bottom_track_149 (
		.in({chanx_right_in[20], bottom_right_grid_left_width_0_height_0_subtile_30__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_37__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_44__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_51__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_58__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_65__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size7_7_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_7_sram_inv[0:2]),
		.out(chany_bottom_out[74]));

	mux_tree_tapbuf_L4SB_size7 mux_bottom_track_163 (
		.in({chanx_right_in[13], bottom_right_grid_left_width_0_height_0_subtile_30__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_37__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_44__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_51__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_58__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_65__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size7_8_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_8_sram_inv[0:2]),
		.out(chany_bottom_out[81]));

	mux_tree_tapbuf_L4SB_size7 mux_bottom_track_177 (
		.in({chanx_right_in[6], bottom_right_grid_left_width_0_height_0_subtile_30__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_37__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_44__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_51__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_58__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_65__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size7_9_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_9_sram_inv[0:2]),
		.out(chany_bottom_out[88]));

	mux_tree_tapbuf_L4SB_size7 mux_bottom_track_191 (
		.in({chanx_right_in[95], bottom_right_grid_left_width_0_height_0_subtile_30__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_37__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_44__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_51__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_58__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_65__pin_a2f_o_0_}),
		.sram(mux_tree_tapbuf_L4SB_size7_10_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_L4SB_size7_10_sram_inv[0:2]),
		.out(chany_bottom_out[95]));

	mux_tree_tapbuf_L4SB_size7_mem mem_bottom_track_51 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size7_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size7_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_0_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7_mem mem_bottom_track_65 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size7_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size7_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_1_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7_mem mem_bottom_track_79 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size7_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size7_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_2_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7_mem mem_bottom_track_93 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size7_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size7_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_3_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7_mem mem_bottom_track_107 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_29_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size7_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size7_4_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_4_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7_mem mem_bottom_track_121 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_35_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size7_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size7_5_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_5_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7_mem mem_bottom_track_135 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_41_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size7_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size7_6_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_6_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7_mem mem_bottom_track_149 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_47_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size7_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size7_7_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_7_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7_mem mem_bottom_track_163 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_53_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size7_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size7_8_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_8_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7_mem mem_bottom_track_177 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_59_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_L4SB_size7_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size7_9_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_9_sram_inv[0:2]));

	mux_tree_tapbuf_L4SB_size7_mem mem_bottom_track_191 (
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.ccff_head(mux_tree_tapbuf_L4SB_size8_mem_65_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mux_tree_tapbuf_L4SB_size7_10_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_L4SB_size7_10_sram_inv[0:2]));

endmodule
// ----- END Verilog module for sb_0__8_ -----

//----- Default net type -----
`default_nettype none



