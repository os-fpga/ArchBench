`default_nettype none

module and8_top_formal_verification_random_tb;

	reg clock0;

	reg [7:0] a;
	wire b;

	wire [0:15] clk;
	wire [0:2303] gfpga_pad_QL_PREIO_A2F;
	wire [0:2303] gfpga_pad_QL_PREIO_F2A;
	wire [0:2303] gfpga_pad_QL_PREIO_F2A_CLK;
	wire [0:513] bl_config_region_0;
	wire [0:406] wl_config_region_0;
	bit global_resetn;
	wire scan_en;
	wire scan_mode;

	fpga_top U0_formal_verification (
		clk[0:15],
		global_resetn,
		scan_en,
		scan_mode,
		gfpga_pad_QL_PREIO_A2F[0:2303],
		gfpga_pad_QL_PREIO_F2A[0:2303],
		gfpga_pad_QL_PREIO_F2A_CLK[0:2303],
		bl_config_region_0[0:513],
		wl_config_region_0[0:406]);

	// assign global_resetn = 1'b0;
	assign scan_en = 1'b0;
	assign scan_mode = 1'b0;
	assign clk[0] = clock0;
	assign clk[1] = 1'b0;
	assign clk[2] = 1'b0;
	assign clk[3] = 1'b0;
	assign clk[4] = 1'b0;
	assign clk[5] = 1'b0;
	assign clk[6] = 1'b0;
	assign clk[7] = 1'b0;
	assign clk[8] = 1'b0;
	assign clk[9] = 1'b0;
	assign clk[10] = 1'b0;
	assign clk[11] = 1'b0;
	assign clk[12] = 1'b0;
	assign clk[13] = 1'b0;
	assign clk[14] = 1'b0;
	assign clk[15] = 1'b0;

	initial begin
		clock0 <= 1'b0;
		while(1) begin
			#1
			clock0 <= !clock0;
		end
	end

	`include "../and8/PinMapping.v"

	initial begin
		`include "../../bitstream_text.txt"
		
		a[0]=1'b0;
		a[1]=1'b0;
		a[2]=1'b0;
		a[3]=1'b0;
		a[4]=1'b0;
		a[5]=1'b0;
		a[6]=1'b0;
		a[7]=1'b0;
		#5;
		global_resetn<=1'b1;
		#5;
		if (b==0)
			$display("Status: Test Passed");
		else
			$display("Status: Test Failed");

		a[0]=1'b1;
		#5;
		if (b==0)
			$display("Status: Test Passed");
		else
			$display("Status: Test Failed");

		a[1]=1'b1;
		#5;
		if (b==0)
			$display("Status: Test Passed");
		else
			$display("Status: Test Failed");

		a[2]=1'b1;
		#5;
		if (b==0)
			$display("Status: Test Passed");
		else
			$display("Status: Test Failed");

		a[3]=1'b1;
		#5;
		if (b==0)
			$display("Status: Test Passed");
		else
			$display("Status: Test Failed");

		a[4]=1'b1;
		#5;
		if (b==0)
			$display("Status: Test Passed");
		else
			$display("Status: Test Failed");

		a[5]=1'b1;
		#5;
		if (b==0)
			$display("Status: Test Passed");
		else
			$display("Status: Test Failed");

		a[6]=1'b1;
		#5;
		if (b==0)
			$display("Status: Test Passed");
		else
			$display("Status: Test Failed");

		a[7]=1'b1;
		#5;
		if (b==1)
			$display("Status: Test Passed");
		else
			$display("Status: Test Failed");
		#10;
		$finish;
	end

	initial begin
		$dumpfile("and8.vcd");
		$dumpvars(1, and8_top_formal_verification_random_tb);
	end

endmodule

