//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for primitive pb_type: logic1
//	Author: Xifan TANG
//	Organization: University of Utah
//-------------------------------------------
//----- Time scale -----
`timescale 1ns / 1ps

//----- Default net type -----
`default_nettype wire

// ----- Verilog module for logical_tile_dsp_mode_default__opt_mode_default__logic1 -----
module logical_tile_dsp_mode_default__opt_mode_default__logic1(logic1_logic1);
//----- OUTPUT PORTS -----
output [0:0] logic1_logic1;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	logic1 logic1_0_ (
		.logic1(logic1_logic1));

endmodule
// ----- END Verilog module for logical_tile_dsp_mode_default__opt_mode_default__logic1 -----

//----- Default net type -----
`default_nettype none



