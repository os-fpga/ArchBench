//--------------------
// Verilog ROM : rom.v
//--------------------
// ROM Specification
//    -8192byte (32bit x 2048word)
//    -module rom(CLK, CE, WE, SEL, ADR, DATI, DATO);
//        input  CLK;         : clock
//        input  CE;          : chip enable
//        input  WE;          : write enable (ignored)
//        input  [ 3:0] SEL;  : byte lane (ignored)
//        input  [12:0] ADR;  : address input
//        input  [31:0] DATI; : data input (ignored)
//        output [31:0] DATO; : data output
//    -CE and ADR are latched at posedge of CLK,
//    -From the negedge of CLK, DAT will be out.
//    -If CE is 0, DAT will be 32'h00000000.
//    -ADR[1:0] are ignored.

`include "../rtl/include/timescale.v"

module rom (CLK, CE, WE, SEL, ADR, DATI, DATO);
    input  CLK, CE, WE;
    input  [ 3:0] SEL;
    input  [12:0] ADR;
    input  [31:0] DATI;
    output [31:0] DATO;

    reg [31:0] DATO;

    always @(negedge CLK) begin
        if (CE == 1'b0)
            DATO <= 32'h00000000;
        else
            begin
                case(ADR[12:2])
                    11'h000 : DATO <= 32'h00000400;
                    11'h001 : DATO <= 32'hFFFD0000;
                    11'h002 : DATO <= 32'h00000000;
                    11'h003 : DATO <= 32'h00000000;
                    11'h004 : DATO <= 32'h00000000;
                    11'h005 : DATO <= 32'h00000000;
                    11'h006 : DATO <= 32'h00000000;
                    11'h007 : DATO <= 32'h00000000;
                    11'h008 : DATO <= 32'h00000000;
                    11'h009 : DATO <= 32'h00000000;
                    11'h00A : DATO <= 32'h00000000;
                    11'h00B : DATO <= 32'h00000000;
                    11'h00C : DATO <= 32'h00000000;
                    11'h00D : DATO <= 32'h00000000;
                    11'h00E : DATO <= 32'h00000000;
                    11'h00F : DATO <= 32'h00000000;
                    11'h010 : DATO <= 32'h00000000;
                    11'h011 : DATO <= 32'h00000000;
                    11'h012 : DATO <= 32'h00000000;
                    11'h013 : DATO <= 32'h00000000;
                    11'h014 : DATO <= 32'h00000000;
                    11'h015 : DATO <= 32'h00000000;
                    11'h016 : DATO <= 32'h00000000;
                    11'h017 : DATO <= 32'h00000000;
                    11'h018 : DATO <= 32'h00000000;
                    11'h019 : DATO <= 32'h00000000;
                    11'h01A : DATO <= 32'h00000000;
                    11'h01B : DATO <= 32'h00000000;
                    11'h01C : DATO <= 32'h00000000;
                    11'h01D : DATO <= 32'h00000000;
                    11'h01E : DATO <= 32'h00000000;
                    11'h01F : DATO <= 32'h00000000;
                    11'h020 : DATO <= 32'h00000000;
                    11'h021 : DATO <= 32'h00000000;
                    11'h022 : DATO <= 32'h00000000;
                    11'h023 : DATO <= 32'h00000000;
                    11'h024 : DATO <= 32'h00000000;
                    11'h025 : DATO <= 32'h00000000;
                    11'h026 : DATO <= 32'h00000000;
                    11'h027 : DATO <= 32'h00000000;
                    11'h028 : DATO <= 32'h00000000;
                    11'h029 : DATO <= 32'h00000000;
                    11'h02A : DATO <= 32'h00000000;
                    11'h02B : DATO <= 32'h00000000;
                    11'h02C : DATO <= 32'h00000000;
                    11'h02D : DATO <= 32'h00000000;
                    11'h02E : DATO <= 32'h00000000;
                    11'h02F : DATO <= 32'h00000000;
                    11'h030 : DATO <= 32'h00000000;
                    11'h031 : DATO <= 32'h00000000;
                    11'h032 : DATO <= 32'h00000000;
                    11'h033 : DATO <= 32'h00000000;
                    11'h034 : DATO <= 32'h00000000;
                    11'h035 : DATO <= 32'h00000000;
                    11'h036 : DATO <= 32'h00000000;
                    11'h037 : DATO <= 32'h00000000;
                    11'h038 : DATO <= 32'h00000000;
                    11'h039 : DATO <= 32'h00000000;
                    11'h03A : DATO <= 32'h00000000;
                    11'h03B : DATO <= 32'h00000000;
                    11'h03C : DATO <= 32'h00000000;
                    11'h03D : DATO <= 32'h00000000;
                    11'h03E : DATO <= 32'h00000000;
                    11'h03F : DATO <= 32'h00000000;
                    11'h040 : DATO <= 32'h00000000;
                    11'h041 : DATO <= 32'h00000000;
                    11'h042 : DATO <= 32'h00000000;
                    11'h043 : DATO <= 32'h00000000;
                    11'h044 : DATO <= 32'h00000000;
                    11'h045 : DATO <= 32'h00000000;
                    11'h046 : DATO <= 32'h00000000;
                    11'h047 : DATO <= 32'h00000000;
                    11'h048 : DATO <= 32'h00000000;
                    11'h049 : DATO <= 32'h00000000;
                    11'h04A : DATO <= 32'h00000000;
                    11'h04B : DATO <= 32'h00000000;
                    11'h04C : DATO <= 32'h00000000;
                    11'h04D : DATO <= 32'h00000000;
                    11'h04E : DATO <= 32'h00000000;
                    11'h04F : DATO <= 32'h00000000;
                    11'h050 : DATO <= 32'h00000000;
                    11'h051 : DATO <= 32'h00000000;
                    11'h052 : DATO <= 32'h00000000;
                    11'h053 : DATO <= 32'h00000000;
                    11'h054 : DATO <= 32'h00000000;
                    11'h055 : DATO <= 32'h00000000;
                    11'h056 : DATO <= 32'h00000000;
                    11'h057 : DATO <= 32'h00000000;
                    11'h058 : DATO <= 32'h00000000;
                    11'h059 : DATO <= 32'h00000000;
                    11'h05A : DATO <= 32'h00000000;
                    11'h05B : DATO <= 32'h00000000;
                    11'h05C : DATO <= 32'h00000000;
                    11'h05D : DATO <= 32'h00000000;
                    11'h05E : DATO <= 32'h00000000;
                    11'h05F : DATO <= 32'h00000000;
                    11'h060 : DATO <= 32'h00000000;
                    11'h061 : DATO <= 32'h00000000;
                    11'h062 : DATO <= 32'h00000000;
                    11'h063 : DATO <= 32'h00000000;
                    11'h064 : DATO <= 32'h00000000;
                    11'h065 : DATO <= 32'h00000000;
                    11'h066 : DATO <= 32'h00000000;
                    11'h067 : DATO <= 32'h00000000;
                    11'h068 : DATO <= 32'h00000000;
                    11'h069 : DATO <= 32'h00000000;
                    11'h06A : DATO <= 32'h00000000;
                    11'h06B : DATO <= 32'h00000000;
                    11'h06C : DATO <= 32'h00000000;
                    11'h06D : DATO <= 32'h00000000;
                    11'h06E : DATO <= 32'h00000000;
                    11'h06F : DATO <= 32'h00000000;
                    11'h070 : DATO <= 32'h00000000;
                    11'h071 : DATO <= 32'h00000000;
                    11'h072 : DATO <= 32'h00000000;
                    11'h073 : DATO <= 32'h00000000;
                    11'h074 : DATO <= 32'h00000000;
                    11'h075 : DATO <= 32'h00000000;
                    11'h076 : DATO <= 32'h00000000;
                    11'h077 : DATO <= 32'h00000000;
                    11'h078 : DATO <= 32'h00000000;
                    11'h079 : DATO <= 32'h00000000;
                    11'h07A : DATO <= 32'h00000000;
                    11'h07B : DATO <= 32'h00000000;
                    11'h07C : DATO <= 32'h00000000;
                    11'h07D : DATO <= 32'h00000000;
                    11'h07E : DATO <= 32'h00000000;
                    11'h07F : DATO <= 32'h00000000;
                    11'h080 : DATO <= 32'h00000000;
                    11'h081 : DATO <= 32'h00000000;
                    11'h082 : DATO <= 32'h00000000;
                    11'h083 : DATO <= 32'h00000000;
                    11'h084 : DATO <= 32'h00000000;
                    11'h085 : DATO <= 32'h00000000;
                    11'h086 : DATO <= 32'h00000000;
                    11'h087 : DATO <= 32'h00000000;
                    11'h088 : DATO <= 32'h00000000;
                    11'h089 : DATO <= 32'h00000000;
                    11'h08A : DATO <= 32'h00000000;
                    11'h08B : DATO <= 32'h00000000;
                    11'h08C : DATO <= 32'h00000000;
                    11'h08D : DATO <= 32'h00000000;
                    11'h08E : DATO <= 32'h00000000;
                    11'h08F : DATO <= 32'h00000000;
                    11'h090 : DATO <= 32'h00000000;
                    11'h091 : DATO <= 32'h00000000;
                    11'h092 : DATO <= 32'h00000000;
                    11'h093 : DATO <= 32'h00000000;
                    11'h094 : DATO <= 32'h00000000;
                    11'h095 : DATO <= 32'h00000000;
                    11'h096 : DATO <= 32'h00000000;
                    11'h097 : DATO <= 32'h00000000;
                    11'h098 : DATO <= 32'h00000000;
                    11'h099 : DATO <= 32'h00000000;
                    11'h09A : DATO <= 32'h00000000;
                    11'h09B : DATO <= 32'h00000000;
                    11'h09C : DATO <= 32'h00000000;
                    11'h09D : DATO <= 32'h00000000;
                    11'h09E : DATO <= 32'h00000000;
                    11'h09F : DATO <= 32'h00000000;
                    11'h0A0 : DATO <= 32'h00000000;
                    11'h0A1 : DATO <= 32'h00000000;
                    11'h0A2 : DATO <= 32'h00000000;
                    11'h0A3 : DATO <= 32'h00000000;
                    11'h0A4 : DATO <= 32'h00000000;
                    11'h0A5 : DATO <= 32'h00000000;
                    11'h0A6 : DATO <= 32'h00000000;
                    11'h0A7 : DATO <= 32'h00000000;
                    11'h0A8 : DATO <= 32'h00000000;
                    11'h0A9 : DATO <= 32'h00000000;
                    11'h0AA : DATO <= 32'h00000000;
                    11'h0AB : DATO <= 32'h00000000;
                    11'h0AC : DATO <= 32'h00000000;
                    11'h0AD : DATO <= 32'h00000000;
                    11'h0AE : DATO <= 32'h00000000;
                    11'h0AF : DATO <= 32'h00000000;
                    11'h0B0 : DATO <= 32'h00000000;
                    11'h0B1 : DATO <= 32'h00000000;
                    11'h0B2 : DATO <= 32'h00000000;
                    11'h0B3 : DATO <= 32'h00000000;
                    11'h0B4 : DATO <= 32'h00000000;
                    11'h0B5 : DATO <= 32'h00000000;
                    11'h0B6 : DATO <= 32'h00000000;
                    11'h0B7 : DATO <= 32'h00000000;
                    11'h0B8 : DATO <= 32'h00000000;
                    11'h0B9 : DATO <= 32'h00000000;
                    11'h0BA : DATO <= 32'h00000000;
                    11'h0BB : DATO <= 32'h00000000;
                    11'h0BC : DATO <= 32'h00000000;
                    11'h0BD : DATO <= 32'h00000000;
                    11'h0BE : DATO <= 32'h00000000;
                    11'h0BF : DATO <= 32'h00000000;
                    11'h0C0 : DATO <= 32'h00000000;
                    11'h0C1 : DATO <= 32'h00000000;
                    11'h0C2 : DATO <= 32'h00000000;
                    11'h0C3 : DATO <= 32'h00000000;
                    11'h0C4 : DATO <= 32'h00000000;
                    11'h0C5 : DATO <= 32'h00000000;
                    11'h0C6 : DATO <= 32'h00000000;
                    11'h0C7 : DATO <= 32'h00000000;
                    11'h0C8 : DATO <= 32'h00000000;
                    11'h0C9 : DATO <= 32'h00000000;
                    11'h0CA : DATO <= 32'h00000000;
                    11'h0CB : DATO <= 32'h00000000;
                    11'h0CC : DATO <= 32'h00000000;
                    11'h0CD : DATO <= 32'h00000000;
                    11'h0CE : DATO <= 32'h00000000;
                    11'h0CF : DATO <= 32'h00000000;
                    11'h0D0 : DATO <= 32'h00000000;
                    11'h0D1 : DATO <= 32'h00000000;
                    11'h0D2 : DATO <= 32'h00000000;
                    11'h0D3 : DATO <= 32'h00000000;
                    11'h0D4 : DATO <= 32'h00000000;
                    11'h0D5 : DATO <= 32'h00000000;
                    11'h0D6 : DATO <= 32'h00000000;
                    11'h0D7 : DATO <= 32'h00000000;
                    11'h0D8 : DATO <= 32'h00000000;
                    11'h0D9 : DATO <= 32'h00000000;
                    11'h0DA : DATO <= 32'h00000000;
                    11'h0DB : DATO <= 32'h00000000;
                    11'h0DC : DATO <= 32'h00000000;
                    11'h0DD : DATO <= 32'h00000000;
                    11'h0DE : DATO <= 32'h00000000;
                    11'h0DF : DATO <= 32'h00000000;
                    11'h0E0 : DATO <= 32'h00000000;
                    11'h0E1 : DATO <= 32'h00000000;
                    11'h0E2 : DATO <= 32'h00000000;
                    11'h0E3 : DATO <= 32'h00000000;
                    11'h0E4 : DATO <= 32'h00000000;
                    11'h0E5 : DATO <= 32'h00000000;
                    11'h0E6 : DATO <= 32'h00000000;
                    11'h0E7 : DATO <= 32'h00000000;
                    11'h0E8 : DATO <= 32'h00000000;
                    11'h0E9 : DATO <= 32'h00000000;
                    11'h0EA : DATO <= 32'h00000000;
                    11'h0EB : DATO <= 32'h00000000;
                    11'h0EC : DATO <= 32'h00000000;
                    11'h0ED : DATO <= 32'h00000000;
                    11'h0EE : DATO <= 32'h00000000;
                    11'h0EF : DATO <= 32'h00000000;
                    11'h0F0 : DATO <= 32'h00000000;
                    11'h0F1 : DATO <= 32'h00000000;
                    11'h0F2 : DATO <= 32'h00000000;
                    11'h0F3 : DATO <= 32'h00000000;
                    11'h0F4 : DATO <= 32'h00000000;
                    11'h0F5 : DATO <= 32'h00000000;
                    11'h0F6 : DATO <= 32'h00000000;
                    11'h0F7 : DATO <= 32'h00000000;
                    11'h0F8 : DATO <= 32'h00000000;
                    11'h0F9 : DATO <= 32'h00000000;
                    11'h0FA : DATO <= 32'h00000000;
                    11'h0FB : DATO <= 32'h00000000;
                    11'h0FC : DATO <= 32'h00000000;
                    11'h0FD : DATO <= 32'h00000000;
                    11'h0FE : DATO <= 32'h00000000;
                    11'h0FF : DATO <= 32'h00000000;
                    11'h100 : DATO <= 32'hEE00DD01;
                    11'h101 : DATO <= 32'hA0020009;
                    11'h102 : DATO <= 32'h00000894;
                    11'h103 : DATO <= 32'hD014620C;
                    11'h104 : DATO <= 32'h640D660E;
                    11'h105 : DATO <= 32'h680FD114;
                    11'h106 : DATO <= 32'hD314D513;
                    11'h107 : DATO <= 32'hD7133210;
                    11'h108 : DATO <= 32'h8B183430;
                    11'h109 : DATO <= 32'h8B163650;
                    11'h10A : DATO <= 32'h8B143870;
                    11'h10B : DATO <= 32'h8B12D00D;
                    11'h10C : DATO <= 32'h620C640D;
                    11'h10D : DATO <= 32'h660E680F;
                    11'h10E : DATO <= 32'hD10DD30E;
                    11'h10F : DATO <= 32'hD50ED70F;
                    11'h110 : DATO <= 32'h32108B07;
                    11'h111 : DATO <= 32'h34308B05;
                    11'h112 : DATO <= 32'h36508B03;
                    11'h113 : DATO <= 32'h38708B01;
                    11'h114 : DATO <= 32'hA0160009;
                    11'h115 : DATO <= 32'h4D2B0009;
                    11'h116 : DATO <= 32'h00090009;
                    11'h117 : DATO <= 32'h00090009;
                    11'h118 : DATO <= 32'h11223344;
                    11'h119 : DATO <= 32'hAABBCCDD;
                    11'h11A : DATO <= 32'h00000044;
                    11'h11B : DATO <= 32'h00003344;
                    11'h11C : DATO <= 32'h000000DD;
                    11'h11D : DATO <= 32'h0000CCDD;
                    11'h11E : DATO <= 32'hFFFFFFDD;
                    11'h11F : DATO <= 32'hFFFFCCDD;
                    11'h120 : DATO <= 32'h0008E400;
                    11'h121 : DATO <= 32'hE201662A;
                    11'h122 : DATO <= 32'h89014D2B;
                    11'h123 : DATO <= 32'h0009684A;
                    11'h124 : DATO <= 32'h89014D2B;
                    11'h125 : DATO <= 32'h0009E4FF;
                    11'h126 : DATO <= 32'hE2FF3480;
                    11'h127 : DATO <= 32'h89014D2B;
                    11'h128 : DATO <= 32'h00093260;
                    11'h129 : DATO <= 32'h89014D2B;
                    11'h12A : DATO <= 32'h00090008;
                    11'h12B : DATO <= 32'hE200602A;
                    11'h12C : DATO <= 32'h8B014D2B;
                    11'h12D : DATO <= 32'h00098800;
                    11'h12E : DATO <= 32'h89014D2B;
                    11'h12F : DATO <= 32'h0009E27F;
                    11'h130 : DATO <= 32'h602B8881;
                    11'h131 : DATO <= 32'h89014D2B;
                    11'h132 : DATO <= 32'h0009E280;
                    11'h133 : DATO <= 32'h602BD404;
                    11'h134 : DATO <= 32'h30408901;
                    11'h135 : DATO <= 32'h4D2B0009;
                    11'h136 : DATO <= 32'hA0040009;
                    11'h137 : DATO <= 32'h00090009;
                    11'h138 : DATO <= 32'h00000080;
                    11'h139 : DATO <= 32'hD2D96428;
                    11'h13A : DATO <= 32'h6629D8DB;
                    11'h13B : DATO <= 32'hDADB3480;
                    11'h13C : DATO <= 32'h89014D2B;
                    11'h13D : DATO <= 32'h000936A0;
                    11'h13E : DATO <= 32'h89014D2B;
                    11'h13F : DATO <= 32'h0009E2AA;
                    11'h140 : DATO <= 32'h60278855;
                    11'h141 : DATO <= 32'h89014D2B;
                    11'h142 : DATO <= 32'h0009D1CD;
                    11'h143 : DATO <= 32'hE0552100;
                    11'h144 : DATO <= 32'h411B8B01;
                    11'h145 : DATO <= 32'h4D2B0009;
                    11'h146 : DATO <= 32'h601088D5;
                    11'h147 : DATO <= 32'h89014D2B;
                    11'h148 : DATO <= 32'h0009E000;
                    11'h149 : DATO <= 32'h2100411B;
                    11'h14A : DATO <= 32'h89014D2B;
                    11'h14B : DATO <= 32'h00096010;
                    11'h14C : DATO <= 32'h88808901;
                    11'h14D : DATO <= 32'h4D2B0009;
                    11'h14E : DATO <= 32'hE200E60A;
                    11'h14F : DATO <= 32'h326C4610;
                    11'h150 : DATO <= 32'h8BFC6023;
                    11'h151 : DATO <= 32'h88378901;
                    11'h152 : DATO <= 32'h4D2B0009;
                    11'h153 : DATO <= 32'hE07EE27F;
                    11'h154 : DATO <= 32'h302B8B01;
                    11'h155 : DATO <= 32'h4D2B0009;
                    11'h156 : DATO <= 32'h88FF8901;
                    11'h157 : DATO <= 32'h4D2B0009;
                    11'h158 : DATO <= 32'hD0B9E201;
                    11'h159 : DATO <= 32'h302B8901;
                    11'h15A : DATO <= 32'h4D2B0009;
                    11'h15B : DATO <= 32'hD2B53020;
                    11'h15C : DATO <= 32'h89014D2B;
                    11'h15D : DATO <= 32'h0009D0B3;
                    11'h15E : DATO <= 32'hE2FF302B;
                    11'h15F : DATO <= 32'h89014D2B;
                    11'h160 : DATO <= 32'h0009D2B1;
                    11'h161 : DATO <= 32'h30208901;
                    11'h162 : DATO <= 32'h4D2B0009;
                    11'h163 : DATO <= 32'h0008E001;
                    11'h164 : DATO <= 32'hE102301A;
                    11'h165 : DATO <= 32'h89014D2B;
                    11'h166 : DATO <= 32'h000988FF;
                    11'h167 : DATO <= 32'h89014D2B;
                    11'h168 : DATO <= 32'h00090018;
                    11'h169 : DATO <= 32'hE004E102;
                    11'h16A : DATO <= 32'h301A8B01;
                    11'h16B : DATO <= 32'h4D2B0009;
                    11'h16C : DATO <= 32'h88018901;
                    11'h16D : DATO <= 32'h4D2B0009;
                    11'h16E : DATO <= 32'hE056E17F;
                    11'h16F : DATO <= 32'h301888D7;
                    11'h170 : DATO <= 32'h89014D2B;
                    11'h171 : DATO <= 32'h0009E012;
                    11'h172 : DATO <= 32'h70348846;
                    11'h173 : DATO <= 32'h89014D2B;
                    11'h174 : DATO <= 32'h00097001;
                    11'h175 : DATO <= 32'h88478901;
                    11'h176 : DATO <= 32'h4D2B0009;
                    11'h177 : DATO <= 32'hE0FFE201;
                    11'h178 : DATO <= 32'h302F8B01;
                    11'h179 : DATO <= 32'h4D2B0009;
                    11'h17A : DATO <= 32'h88008901;
                    11'h17B : DATO <= 32'h4D2B0009;
                    11'h17C : DATO <= 32'hD094E201;
                    11'h17D : DATO <= 32'h302F8901;
                    11'h17E : DATO <= 32'h4D2B0009;
                    11'h17F : DATO <= 32'hD2923020;
                    11'h180 : DATO <= 32'h89014D2B;
                    11'h181 : DATO <= 32'h0009D090;
                    11'h182 : DATO <= 32'hE2FF302F;
                    11'h183 : DATO <= 32'h89014D2B;
                    11'h184 : DATO <= 32'h0009D28C;
                    11'h185 : DATO <= 32'h30208901;
                    11'h186 : DATO <= 32'h4D2B0009;
                    11'h187 : DATO <= 32'h0008E0FF;
                    11'h188 : DATO <= 32'hE101301E;
                    11'h189 : DATO <= 32'h89014D2B;
                    11'h18A : DATO <= 32'h00098800;
                    11'h18B : DATO <= 32'h89014D2B;
                    11'h18C : DATO <= 32'h00090018;
                    11'h18D : DATO <= 32'hE0FDE101;
                    11'h18E : DATO <= 32'h301E8B01;
                    11'h18F : DATO <= 32'h4D2B0009;
                    11'h190 : DATO <= 32'h88FF8901;
                    11'h191 : DATO <= 32'h4D2B0009;
                    11'h192 : DATO <= 32'hE059E180;
                    11'h193 : DATO <= 32'h301C88D9;
                    11'h194 : DATO <= 32'h89014D2B;
                    11'h195 : DATO <= 32'h0009D27D;
                    11'h196 : DATO <= 32'hD47D224D;
                    11'h197 : DATO <= 32'hD67D3260;
                    11'h198 : DATO <= 32'h89014D2B;
                    11'h199 : DATO <= 32'h0009E0AA;
                    11'h19A : DATO <= 32'hE255202A;
                    11'h19B : DATO <= 32'hC8008901;
                    11'h19C : DATO <= 32'h4D2B0009;
                    11'h19D : DATO <= 32'hE0AAE277;
                    11'h19E : DATO <= 32'h202A88DD;
                    11'h19F : DATO <= 32'h89014D2B;
                    11'h1A0 : DATO <= 32'h0009D16F;
                    11'h1A1 : DATO <= 32'h411EE0AA;
                    11'h1A2 : DATO <= 32'h8017E007;
                    11'h1A3 : DATO <= 32'hCE558417;
                    11'h1A4 : DATO <= 32'h88FF8901;
                    11'h1A5 : DATO <= 32'h4D2B0009;
                    11'h1A6 : DATO <= 32'hE0AA8017;
                    11'h1A7 : DATO <= 32'hE007CE77;
                    11'h1A8 : DATO <= 32'h841788DD;
                    11'h1A9 : DATO <= 32'h89014D2B;
                    11'h1AA : DATO <= 32'h0009E2AA;
                    11'h1AB : DATO <= 32'hE4552248;
                    11'h1AC : DATO <= 32'h00298801;
                    11'h1AD : DATO <= 32'h89014D2B;
                    11'h1AE : DATO <= 32'h0009E2AA;
                    11'h1AF : DATO <= 32'hE45D2248;
                    11'h1B0 : DATO <= 32'h00298800;
                    11'h1B1 : DATO <= 32'h89014D2B;
                    11'h1B2 : DATO <= 32'h0009E0AA;
                    11'h1B3 : DATO <= 32'hC8550029;
                    11'h1B4 : DATO <= 32'h88018901;
                    11'h1B5 : DATO <= 32'h4D2B0009;
                    11'h1B6 : DATO <= 32'hE0AAC8D5;
                    11'h1B7 : DATO <= 32'h00298800;
                    11'h1B8 : DATO <= 32'h89014D2B;
                    11'h1B9 : DATO <= 32'h0009D156;
                    11'h1BA : DATO <= 32'h411EE0AA;
                    11'h1BB : DATO <= 32'h8019E009;
                    11'h1BC : DATO <= 32'h0008CC55;
                    11'h1BD : DATO <= 32'h89014D2B;
                    11'h1BE : DATO <= 32'h0009E0AA;
                    11'h1BF : DATO <= 32'h801BE00B;
                    11'h1C0 : DATO <= 32'h0018CCD5;
                    11'h1C1 : DATO <= 32'h8B014D2B;
                    11'h1C2 : DATO <= 32'h0009E000;
                    11'h1C3 : DATO <= 32'hE1FF2019;
                    11'h1C4 : DATO <= 32'h88008901;
                    11'h1C5 : DATO <= 32'h4D2B0009;
                    11'h1C6 : DATO <= 32'hE0AAE155;
                    11'h1C7 : DATO <= 32'h20198800;
                    11'h1C8 : DATO <= 32'h89014D2B;
                    11'h1C9 : DATO <= 32'h0009E07E;
                    11'h1CA : DATO <= 32'hE1DB2019;
                    11'h1CB : DATO <= 32'h885A8901;
                    11'h1CC : DATO <= 32'h4D2B0009;
                    11'h1CD : DATO <= 32'hE000C9FF;
                    11'h1CE : DATO <= 32'h88008901;
                    11'h1CF : DATO <= 32'h4D2B0009;
                    11'h1D0 : DATO <= 32'hE0AAC955;
                    11'h1D1 : DATO <= 32'h88008901;
                    11'h1D2 : DATO <= 32'h4D2B0009;
                    11'h1D3 : DATO <= 32'hE07EC9DB;
                    11'h1D4 : DATO <= 32'h885A8901;
                    11'h1D5 : DATO <= 32'h4D2B0009;
                    11'h1D6 : DATO <= 32'hD139411E;
                    11'h1D7 : DATO <= 32'hE0008017;
                    11'h1D8 : DATO <= 32'hE007CDFF;
                    11'h1D9 : DATO <= 32'h84178800;
                    11'h1DA : DATO <= 32'h89014D2B;
                    11'h1DB : DATO <= 32'h0009E0AA;
                    11'h1DC : DATO <= 32'h8017E007;
                    11'h1DD : DATO <= 32'hCD558417;
                    11'h1DE : DATO <= 32'h88008901;
                    11'h1DF : DATO <= 32'h4D2B0009;
                    11'h1E0 : DATO <= 32'hE07E8017;
                    11'h1E1 : DATO <= 32'hE007CDDB;
                    11'h1E2 : DATO <= 32'h8417885A;
                    11'h1E3 : DATO <= 32'h89014D2B;
                    11'h1E4 : DATO <= 32'h0009E000;
                    11'h1E5 : DATO <= 32'hE1FF201B;
                    11'h1E6 : DATO <= 32'h88FF8901;
                    11'h1E7 : DATO <= 32'h4D2B0009;
                    11'h1E8 : DATO <= 32'hE0AAE155;
                    11'h1E9 : DATO <= 32'h201B88FF;
                    11'h1EA : DATO <= 32'h89014D2B;
                    11'h1EB : DATO <= 32'h0009E055;
                    11'h1EC : DATO <= 32'hE15A201B;
                    11'h1ED : DATO <= 32'h885F8901;
                    11'h1EE : DATO <= 32'h4D2B0009;
                    11'h1EF : DATO <= 32'hE000CBFF;
                    11'h1F0 : DATO <= 32'h924E3020;
                    11'h1F1 : DATO <= 32'h89014D2B;
                    11'h1F2 : DATO <= 32'h0009E0AA;
                    11'h1F3 : DATO <= 32'hCB559248;
                    11'h1F4 : DATO <= 32'h30208901;
                    11'h1F5 : DATO <= 32'h4D2B0009;
                    11'h1F6 : DATO <= 32'hE055CB5A;
                    11'h1F7 : DATO <= 32'h885F8901;
                    11'h1F8 : DATO <= 32'h4D2B0009;
                    11'h1F9 : DATO <= 32'hD116411E;
                    11'h1FA : DATO <= 32'hE0008017;
                    11'h1FB : DATO <= 32'hE007CFFF;
                    11'h1FC : DATO <= 32'h841788FF;
                    11'h1FD : DATO <= 32'h89014D2B;
                    11'h1FE : DATO <= 32'h0009E0AA;
                    11'h1FF : DATO <= 32'h8017E007;
                    11'h200 : DATO <= 32'hCF558417;
                    11'h201 : DATO <= 32'h88FF8901;
                    11'h202 : DATO <= 32'h4D2B0009;
                    11'h203 : DATO <= 32'hE0558017;
                    11'h204 : DATO <= 32'hE007CF5A;
                    11'h205 : DATO <= 32'h8417885F;
                    11'h206 : DATO <= 32'h89014D2B;
                    11'h207 : DATO <= 32'h00090018;
                    11'h208 : DATO <= 32'h00298801;
                    11'h209 : DATO <= 32'h89014D2B;
                    11'h20A : DATO <= 32'h00090008;
                    11'h20B : DATO <= 32'h00298800;
                    11'h20C : DATO <= 32'h89014D2B;
                    11'h20D : DATO <= 32'h0009A015;
                    11'h20E : DATO <= 32'h00090009;
                    11'h20F : DATO <= 32'h00090009;
                    11'h210 : DATO <= 32'hFFFCE000;
                    11'h211 : DATO <= 32'h7FFFFFFF;
                    11'h212 : DATO <= 32'h80000000;
                    11'h213 : DATO <= 32'h00112233;
                    11'h214 : DATO <= 32'h44556677;
                    11'h215 : DATO <= 32'h66770011;
                    11'h216 : DATO <= 32'h00113322;
                    11'h217 : DATO <= 32'h22330011;
                    11'h218 : DATO <= 32'h00FFFFFF;
                    11'h219 : DATO <= 32'hDD023DEC;
                    11'h21A : DATO <= 32'h6CD24C2B;
                    11'h21B : DATO <= 32'h7E040009;
                    11'h21C : DATO <= 32'h00000874;
                    11'h21D : DATO <= 32'h00010402;
                    11'h21E : DATO <= 32'h00020402;
                    11'h21F : DATO <= 32'h00030402;
                    11'h220 : DATO <= 32'h00000884;
                    11'h221 : DATO <= 32'hD002D102;
                    11'h222 : DATO <= 32'h2102AFFB;
                    11'h223 : DATO <= 32'h00090009;
                    11'h224 : DATO <= 32'h12345678;
                    11'h225 : DATO <= 32'hD002D102;
                    11'h226 : DATO <= 32'hAFFC0009;
                    11'h227 : DATO <= 32'h00090009;
                    11'h228 : DATO <= 32'h88888888;
                    11'h229 : DATO <= 32'h00090009;
                    11'h22A : DATO <= 32'h00090009;
                    11'h22B : DATO <= 32'h00090009;
                    11'h22C : DATO <= 32'hFFFFFFFF;
                    11'h22D : DATO <= 32'hFFFFFFFF;
                    11'h22E : DATO <= 32'hFFFFFFFF;
                    11'h22F : DATO <= 32'hFFFFFFFF;
                    11'h230 : DATO <= 32'hFFFFFFFF;
                    11'h231 : DATO <= 32'hFFFFFFFF;
                    11'h232 : DATO <= 32'hFFFFFFFF;
                    11'h233 : DATO <= 32'hFFFFFFFF;
                    11'h234 : DATO <= 32'hFFFFFFFF;
                    11'h235 : DATO <= 32'hFFFFFFFF;
                    11'h236 : DATO <= 32'hFFFFFFFF;
                    11'h237 : DATO <= 32'hFFFFFFFF;
                    11'h238 : DATO <= 32'hFFFFFFFF;
                    11'h239 : DATO <= 32'hFFFFFFFF;
                    11'h23A : DATO <= 32'hFFFFFFFF;
                    11'h23B : DATO <= 32'hFFFFFFFF;
                    11'h23C : DATO <= 32'hFFFFFFFF;
                    11'h23D : DATO <= 32'hFFFFFFFF;
                    11'h23E : DATO <= 32'hFFFFFFFF;
                    11'h23F : DATO <= 32'hFFFFFFFF;
                    11'h240 : DATO <= 32'hFFFFFFFF;
                    11'h241 : DATO <= 32'hFFFFFFFF;
                    11'h242 : DATO <= 32'hFFFFFFFF;
                    11'h243 : DATO <= 32'hFFFFFFFF;
                    11'h244 : DATO <= 32'hFFFFFFFF;
                    11'h245 : DATO <= 32'hFFFFFFFF;
                    11'h246 : DATO <= 32'hFFFFFFFF;
                    11'h247 : DATO <= 32'hFFFFFFFF;
                    11'h248 : DATO <= 32'hFFFFFFFF;
                    11'h249 : DATO <= 32'hFFFFFFFF;
                    11'h24A : DATO <= 32'hFFFFFFFF;
                    11'h24B : DATO <= 32'hFFFFFFFF;
                    11'h24C : DATO <= 32'hFFFFFFFF;
                    11'h24D : DATO <= 32'hFFFFFFFF;
                    11'h24E : DATO <= 32'hFFFFFFFF;
                    11'h24F : DATO <= 32'hFFFFFFFF;
                    11'h250 : DATO <= 32'hFFFFFFFF;
                    11'h251 : DATO <= 32'hFFFFFFFF;
                    11'h252 : DATO <= 32'hFFFFFFFF;
                    11'h253 : DATO <= 32'hFFFFFFFF;
                    11'h254 : DATO <= 32'hFFFFFFFF;
                    11'h255 : DATO <= 32'hFFFFFFFF;
                    11'h256 : DATO <= 32'hFFFFFFFF;
                    11'h257 : DATO <= 32'hFFFFFFFF;
                    11'h258 : DATO <= 32'hFFFFFFFF;
                    11'h259 : DATO <= 32'hFFFFFFFF;
                    11'h25A : DATO <= 32'hFFFFFFFF;
                    11'h25B : DATO <= 32'hFFFFFFFF;
                    11'h25C : DATO <= 32'hFFFFFFFF;
                    11'h25D : DATO <= 32'hFFFFFFFF;
                    11'h25E : DATO <= 32'hFFFFFFFF;
                    11'h25F : DATO <= 32'hFFFFFFFF;
                    11'h260 : DATO <= 32'hFFFFFFFF;
                    11'h261 : DATO <= 32'hFFFFFFFF;
                    11'h262 : DATO <= 32'hFFFFFFFF;
                    11'h263 : DATO <= 32'hFFFFFFFF;
                    11'h264 : DATO <= 32'hFFFFFFFF;
                    11'h265 : DATO <= 32'hFFFFFFFF;
                    11'h266 : DATO <= 32'hFFFFFFFF;
                    11'h267 : DATO <= 32'hFFFFFFFF;
                    11'h268 : DATO <= 32'hFFFFFFFF;
                    11'h269 : DATO <= 32'hFFFFFFFF;
                    11'h26A : DATO <= 32'hFFFFFFFF;
                    11'h26B : DATO <= 32'hFFFFFFFF;
                    11'h26C : DATO <= 32'hFFFFFFFF;
                    11'h26D : DATO <= 32'hFFFFFFFF;
                    11'h26E : DATO <= 32'hFFFFFFFF;
                    11'h26F : DATO <= 32'hFFFFFFFF;
                    11'h270 : DATO <= 32'hFFFFFFFF;
                    11'h271 : DATO <= 32'hFFFFFFFF;
                    11'h272 : DATO <= 32'hFFFFFFFF;
                    11'h273 : DATO <= 32'hFFFFFFFF;
                    11'h274 : DATO <= 32'hFFFFFFFF;
                    11'h275 : DATO <= 32'hFFFFFFFF;
                    11'h276 : DATO <= 32'hFFFFFFFF;
                    11'h277 : DATO <= 32'hFFFFFFFF;
                    11'h278 : DATO <= 32'hFFFFFFFF;
                    11'h279 : DATO <= 32'hFFFFFFFF;
                    11'h27A : DATO <= 32'hFFFFFFFF;
                    11'h27B : DATO <= 32'hFFFFFFFF;
                    11'h27C : DATO <= 32'hFFFFFFFF;
                    11'h27D : DATO <= 32'hFFFFFFFF;
                    11'h27E : DATO <= 32'hFFFFFFFF;
                    11'h27F : DATO <= 32'hFFFFFFFF;
                    11'h280 : DATO <= 32'hFFFFFFFF;
                    11'h281 : DATO <= 32'hFFFFFFFF;
                    11'h282 : DATO <= 32'hFFFFFFFF;
                    11'h283 : DATO <= 32'hFFFFFFFF;
                    11'h284 : DATO <= 32'hFFFFFFFF;
                    11'h285 : DATO <= 32'hFFFFFFFF;
                    11'h286 : DATO <= 32'hFFFFFFFF;
                    11'h287 : DATO <= 32'hFFFFFFFF;
                    11'h288 : DATO <= 32'hFFFFFFFF;
                    11'h289 : DATO <= 32'hFFFFFFFF;
                    11'h28A : DATO <= 32'hFFFFFFFF;
                    11'h28B : DATO <= 32'hFFFFFFFF;
                    11'h28C : DATO <= 32'hFFFFFFFF;
                    11'h28D : DATO <= 32'hFFFFFFFF;
                    11'h28E : DATO <= 32'hFFFFFFFF;
                    11'h28F : DATO <= 32'hFFFFFFFF;
                    11'h290 : DATO <= 32'hFFFFFFFF;
                    11'h291 : DATO <= 32'hFFFFFFFF;
                    11'h292 : DATO <= 32'hFFFFFFFF;
                    11'h293 : DATO <= 32'hFFFFFFFF;
                    11'h294 : DATO <= 32'hFFFFFFFF;
                    11'h295 : DATO <= 32'hFFFFFFFF;
                    11'h296 : DATO <= 32'hFFFFFFFF;
                    11'h297 : DATO <= 32'hFFFFFFFF;
                    11'h298 : DATO <= 32'hFFFFFFFF;
                    11'h299 : DATO <= 32'hFFFFFFFF;
                    11'h29A : DATO <= 32'hFFFFFFFF;
                    11'h29B : DATO <= 32'hFFFFFFFF;
                    11'h29C : DATO <= 32'hFFFFFFFF;
                    11'h29D : DATO <= 32'hFFFFFFFF;
                    11'h29E : DATO <= 32'hFFFFFFFF;
                    11'h29F : DATO <= 32'hFFFFFFFF;
                    11'h2A0 : DATO <= 32'hFFFFFFFF;
                    11'h2A1 : DATO <= 32'hFFFFFFFF;
                    11'h2A2 : DATO <= 32'hFFFFFFFF;
                    11'h2A3 : DATO <= 32'hFFFFFFFF;
                    11'h2A4 : DATO <= 32'hFFFFFFFF;
                    11'h2A5 : DATO <= 32'hFFFFFFFF;
                    11'h2A6 : DATO <= 32'hFFFFFFFF;
                    11'h2A7 : DATO <= 32'hFFFFFFFF;
                    11'h2A8 : DATO <= 32'hFFFFFFFF;
                    11'h2A9 : DATO <= 32'hFFFFFFFF;
                    11'h2AA : DATO <= 32'hFFFFFFFF;
                    11'h2AB : DATO <= 32'hFFFFFFFF;
                    11'h2AC : DATO <= 32'hFFFFFFFF;
                    11'h2AD : DATO <= 32'hFFFFFFFF;
                    11'h2AE : DATO <= 32'hFFFFFFFF;
                    11'h2AF : DATO <= 32'hFFFFFFFF;
                    11'h2B0 : DATO <= 32'hFFFFFFFF;
                    11'h2B1 : DATO <= 32'hFFFFFFFF;
                    11'h2B2 : DATO <= 32'hFFFFFFFF;
                    11'h2B3 : DATO <= 32'hFFFFFFFF;
                    11'h2B4 : DATO <= 32'hFFFFFFFF;
                    11'h2B5 : DATO <= 32'hFFFFFFFF;
                    11'h2B6 : DATO <= 32'hFFFFFFFF;
                    11'h2B7 : DATO <= 32'hFFFFFFFF;
                    11'h2B8 : DATO <= 32'hFFFFFFFF;
                    11'h2B9 : DATO <= 32'hFFFFFFFF;
                    11'h2BA : DATO <= 32'hFFFFFFFF;
                    11'h2BB : DATO <= 32'hFFFFFFFF;
                    11'h2BC : DATO <= 32'hFFFFFFFF;
                    11'h2BD : DATO <= 32'hFFFFFFFF;
                    11'h2BE : DATO <= 32'hFFFFFFFF;
                    11'h2BF : DATO <= 32'hFFFFFFFF;
                    11'h2C0 : DATO <= 32'hFFFFFFFF;
                    11'h2C1 : DATO <= 32'hFFFFFFFF;
                    11'h2C2 : DATO <= 32'hFFFFFFFF;
                    11'h2C3 : DATO <= 32'hFFFFFFFF;
                    11'h2C4 : DATO <= 32'hFFFFFFFF;
                    11'h2C5 : DATO <= 32'hFFFFFFFF;
                    11'h2C6 : DATO <= 32'hFFFFFFFF;
                    11'h2C7 : DATO <= 32'hFFFFFFFF;
                    11'h2C8 : DATO <= 32'hFFFFFFFF;
                    11'h2C9 : DATO <= 32'hFFFFFFFF;
                    11'h2CA : DATO <= 32'hFFFFFFFF;
                    11'h2CB : DATO <= 32'hFFFFFFFF;
                    11'h2CC : DATO <= 32'hFFFFFFFF;
                    11'h2CD : DATO <= 32'hFFFFFFFF;
                    11'h2CE : DATO <= 32'hFFFFFFFF;
                    11'h2CF : DATO <= 32'hFFFFFFFF;
                    11'h2D0 : DATO <= 32'hFFFFFFFF;
                    11'h2D1 : DATO <= 32'hFFFFFFFF;
                    11'h2D2 : DATO <= 32'hFFFFFFFF;
                    11'h2D3 : DATO <= 32'hFFFFFFFF;
                    11'h2D4 : DATO <= 32'hFFFFFFFF;
                    11'h2D5 : DATO <= 32'hFFFFFFFF;
                    11'h2D6 : DATO <= 32'hFFFFFFFF;
                    11'h2D7 : DATO <= 32'hFFFFFFFF;
                    11'h2D8 : DATO <= 32'hFFFFFFFF;
                    11'h2D9 : DATO <= 32'hFFFFFFFF;
                    11'h2DA : DATO <= 32'hFFFFFFFF;
                    11'h2DB : DATO <= 32'hFFFFFFFF;
                    11'h2DC : DATO <= 32'hFFFFFFFF;
                    11'h2DD : DATO <= 32'hFFFFFFFF;
                    11'h2DE : DATO <= 32'hFFFFFFFF;
                    11'h2DF : DATO <= 32'hFFFFFFFF;
                    11'h2E0 : DATO <= 32'hFFFFFFFF;
                    11'h2E1 : DATO <= 32'hFFFFFFFF;
                    11'h2E2 : DATO <= 32'hFFFFFFFF;
                    11'h2E3 : DATO <= 32'hFFFFFFFF;
                    11'h2E4 : DATO <= 32'hFFFFFFFF;
                    11'h2E5 : DATO <= 32'hFFFFFFFF;
                    11'h2E6 : DATO <= 32'hFFFFFFFF;
                    11'h2E7 : DATO <= 32'hFFFFFFFF;
                    11'h2E8 : DATO <= 32'hFFFFFFFF;
                    11'h2E9 : DATO <= 32'hFFFFFFFF;
                    11'h2EA : DATO <= 32'hFFFFFFFF;
                    11'h2EB : DATO <= 32'hFFFFFFFF;
                    11'h2EC : DATO <= 32'hFFFFFFFF;
                    11'h2ED : DATO <= 32'hFFFFFFFF;
                    11'h2EE : DATO <= 32'hFFFFFFFF;
                    11'h2EF : DATO <= 32'hFFFFFFFF;
                    11'h2F0 : DATO <= 32'hFFFFFFFF;
                    11'h2F1 : DATO <= 32'hFFFFFFFF;
                    11'h2F2 : DATO <= 32'hFFFFFFFF;
                    11'h2F3 : DATO <= 32'hFFFFFFFF;
                    11'h2F4 : DATO <= 32'hFFFFFFFF;
                    11'h2F5 : DATO <= 32'hFFFFFFFF;
                    11'h2F6 : DATO <= 32'hFFFFFFFF;
                    11'h2F7 : DATO <= 32'hFFFFFFFF;
                    11'h2F8 : DATO <= 32'hFFFFFFFF;
                    11'h2F9 : DATO <= 32'hFFFFFFFF;
                    11'h2FA : DATO <= 32'hFFFFFFFF;
                    11'h2FB : DATO <= 32'hFFFFFFFF;
                    11'h2FC : DATO <= 32'hFFFFFFFF;
                    11'h2FD : DATO <= 32'hFFFFFFFF;
                    11'h2FE : DATO <= 32'hFFFFFFFF;
                    11'h2FF : DATO <= 32'hFFFFFFFF;
                    11'h300 : DATO <= 32'hFFFFFFFF;
                    11'h301 : DATO <= 32'hFFFFFFFF;
                    11'h302 : DATO <= 32'hFFFFFFFF;
                    11'h303 : DATO <= 32'hFFFFFFFF;
                    11'h304 : DATO <= 32'hFFFFFFFF;
                    11'h305 : DATO <= 32'hFFFFFFFF;
                    11'h306 : DATO <= 32'hFFFFFFFF;
                    11'h307 : DATO <= 32'hFFFFFFFF;
                    11'h308 : DATO <= 32'hFFFFFFFF;
                    11'h309 : DATO <= 32'hFFFFFFFF;
                    11'h30A : DATO <= 32'hFFFFFFFF;
                    11'h30B : DATO <= 32'hFFFFFFFF;
                    11'h30C : DATO <= 32'hFFFFFFFF;
                    11'h30D : DATO <= 32'hFFFFFFFF;
                    11'h30E : DATO <= 32'hFFFFFFFF;
                    11'h30F : DATO <= 32'hFFFFFFFF;
                    11'h310 : DATO <= 32'hFFFFFFFF;
                    11'h311 : DATO <= 32'hFFFFFFFF;
                    11'h312 : DATO <= 32'hFFFFFFFF;
                    11'h313 : DATO <= 32'hFFFFFFFF;
                    11'h314 : DATO <= 32'hFFFFFFFF;
                    11'h315 : DATO <= 32'hFFFFFFFF;
                    11'h316 : DATO <= 32'hFFFFFFFF;
                    11'h317 : DATO <= 32'hFFFFFFFF;
                    11'h318 : DATO <= 32'hFFFFFFFF;
                    11'h319 : DATO <= 32'hFFFFFFFF;
                    11'h31A : DATO <= 32'hFFFFFFFF;
                    11'h31B : DATO <= 32'hFFFFFFFF;
                    11'h31C : DATO <= 32'hFFFFFFFF;
                    11'h31D : DATO <= 32'hFFFFFFFF;
                    11'h31E : DATO <= 32'hFFFFFFFF;
                    11'h31F : DATO <= 32'hFFFFFFFF;
                    11'h320 : DATO <= 32'hFFFFFFFF;
                    11'h321 : DATO <= 32'hFFFFFFFF;
                    11'h322 : DATO <= 32'hFFFFFFFF;
                    11'h323 : DATO <= 32'hFFFFFFFF;
                    11'h324 : DATO <= 32'hFFFFFFFF;
                    11'h325 : DATO <= 32'hFFFFFFFF;
                    11'h326 : DATO <= 32'hFFFFFFFF;
                    11'h327 : DATO <= 32'hFFFFFFFF;
                    11'h328 : DATO <= 32'hFFFFFFFF;
                    11'h329 : DATO <= 32'hFFFFFFFF;
                    11'h32A : DATO <= 32'hFFFFFFFF;
                    11'h32B : DATO <= 32'hFFFFFFFF;
                    11'h32C : DATO <= 32'hFFFFFFFF;
                    11'h32D : DATO <= 32'hFFFFFFFF;
                    11'h32E : DATO <= 32'hFFFFFFFF;
                    11'h32F : DATO <= 32'hFFFFFFFF;
                    11'h330 : DATO <= 32'hFFFFFFFF;
                    11'h331 : DATO <= 32'hFFFFFFFF;
                    11'h332 : DATO <= 32'hFFFFFFFF;
                    11'h333 : DATO <= 32'hFFFFFFFF;
                    11'h334 : DATO <= 32'hFFFFFFFF;
                    11'h335 : DATO <= 32'hFFFFFFFF;
                    11'h336 : DATO <= 32'hFFFFFFFF;
                    11'h337 : DATO <= 32'hFFFFFFFF;
                    11'h338 : DATO <= 32'hFFFFFFFF;
                    11'h339 : DATO <= 32'hFFFFFFFF;
                    11'h33A : DATO <= 32'hFFFFFFFF;
                    11'h33B : DATO <= 32'hFFFFFFFF;
                    11'h33C : DATO <= 32'hFFFFFFFF;
                    11'h33D : DATO <= 32'hFFFFFFFF;
                    11'h33E : DATO <= 32'hFFFFFFFF;
                    11'h33F : DATO <= 32'hFFFFFFFF;
                    11'h340 : DATO <= 32'hFFFFFFFF;
                    11'h341 : DATO <= 32'hFFFFFFFF;
                    11'h342 : DATO <= 32'hFFFFFFFF;
                    11'h343 : DATO <= 32'hFFFFFFFF;
                    11'h344 : DATO <= 32'hFFFFFFFF;
                    11'h345 : DATO <= 32'hFFFFFFFF;
                    11'h346 : DATO <= 32'hFFFFFFFF;
                    11'h347 : DATO <= 32'hFFFFFFFF;
                    11'h348 : DATO <= 32'hFFFFFFFF;
                    11'h349 : DATO <= 32'hFFFFFFFF;
                    11'h34A : DATO <= 32'hFFFFFFFF;
                    11'h34B : DATO <= 32'hFFFFFFFF;
                    11'h34C : DATO <= 32'hFFFFFFFF;
                    11'h34D : DATO <= 32'hFFFFFFFF;
                    11'h34E : DATO <= 32'hFFFFFFFF;
                    11'h34F : DATO <= 32'hFFFFFFFF;
                    11'h350 : DATO <= 32'hFFFFFFFF;
                    11'h351 : DATO <= 32'hFFFFFFFF;
                    11'h352 : DATO <= 32'hFFFFFFFF;
                    11'h353 : DATO <= 32'hFFFFFFFF;
                    11'h354 : DATO <= 32'hFFFFFFFF;
                    11'h355 : DATO <= 32'hFFFFFFFF;
                    11'h356 : DATO <= 32'hFFFFFFFF;
                    11'h357 : DATO <= 32'hFFFFFFFF;
                    11'h358 : DATO <= 32'hFFFFFFFF;
                    11'h359 : DATO <= 32'hFFFFFFFF;
                    11'h35A : DATO <= 32'hFFFFFFFF;
                    11'h35B : DATO <= 32'hFFFFFFFF;
                    11'h35C : DATO <= 32'hFFFFFFFF;
                    11'h35D : DATO <= 32'hFFFFFFFF;
                    11'h35E : DATO <= 32'hFFFFFFFF;
                    11'h35F : DATO <= 32'hFFFFFFFF;
                    11'h360 : DATO <= 32'hFFFFFFFF;
                    11'h361 : DATO <= 32'hFFFFFFFF;
                    11'h362 : DATO <= 32'hFFFFFFFF;
                    11'h363 : DATO <= 32'hFFFFFFFF;
                    11'h364 : DATO <= 32'hFFFFFFFF;
                    11'h365 : DATO <= 32'hFFFFFFFF;
                    11'h366 : DATO <= 32'hFFFFFFFF;
                    11'h367 : DATO <= 32'hFFFFFFFF;
                    11'h368 : DATO <= 32'hFFFFFFFF;
                    11'h369 : DATO <= 32'hFFFFFFFF;
                    11'h36A : DATO <= 32'hFFFFFFFF;
                    11'h36B : DATO <= 32'hFFFFFFFF;
                    11'h36C : DATO <= 32'hFFFFFFFF;
                    11'h36D : DATO <= 32'hFFFFFFFF;
                    11'h36E : DATO <= 32'hFFFFFFFF;
                    11'h36F : DATO <= 32'hFFFFFFFF;
                    11'h370 : DATO <= 32'hFFFFFFFF;
                    11'h371 : DATO <= 32'hFFFFFFFF;
                    11'h372 : DATO <= 32'hFFFFFFFF;
                    11'h373 : DATO <= 32'hFFFFFFFF;
                    11'h374 : DATO <= 32'hFFFFFFFF;
                    11'h375 : DATO <= 32'hFFFFFFFF;
                    11'h376 : DATO <= 32'hFFFFFFFF;
                    11'h377 : DATO <= 32'hFFFFFFFF;
                    11'h378 : DATO <= 32'hFFFFFFFF;
                    11'h379 : DATO <= 32'hFFFFFFFF;
                    11'h37A : DATO <= 32'hFFFFFFFF;
                    11'h37B : DATO <= 32'hFFFFFFFF;
                    11'h37C : DATO <= 32'hFFFFFFFF;
                    11'h37D : DATO <= 32'hFFFFFFFF;
                    11'h37E : DATO <= 32'hFFFFFFFF;
                    11'h37F : DATO <= 32'hFFFFFFFF;
                    11'h380 : DATO <= 32'hFFFFFFFF;
                    11'h381 : DATO <= 32'hFFFFFFFF;
                    11'h382 : DATO <= 32'hFFFFFFFF;
                    11'h383 : DATO <= 32'hFFFFFFFF;
                    11'h384 : DATO <= 32'hFFFFFFFF;
                    11'h385 : DATO <= 32'hFFFFFFFF;
                    11'h386 : DATO <= 32'hFFFFFFFF;
                    11'h387 : DATO <= 32'hFFFFFFFF;
                    11'h388 : DATO <= 32'hFFFFFFFF;
                    11'h389 : DATO <= 32'hFFFFFFFF;
                    11'h38A : DATO <= 32'hFFFFFFFF;
                    11'h38B : DATO <= 32'hFFFFFFFF;
                    11'h38C : DATO <= 32'hFFFFFFFF;
                    11'h38D : DATO <= 32'hFFFFFFFF;
                    11'h38E : DATO <= 32'hFFFFFFFF;
                    11'h38F : DATO <= 32'hFFFFFFFF;
                    11'h390 : DATO <= 32'hFFFFFFFF;
                    11'h391 : DATO <= 32'hFFFFFFFF;
                    11'h392 : DATO <= 32'hFFFFFFFF;
                    11'h393 : DATO <= 32'hFFFFFFFF;
                    11'h394 : DATO <= 32'hFFFFFFFF;
                    11'h395 : DATO <= 32'hFFFFFFFF;
                    11'h396 : DATO <= 32'hFFFFFFFF;
                    11'h397 : DATO <= 32'hFFFFFFFF;
                    11'h398 : DATO <= 32'hFFFFFFFF;
                    11'h399 : DATO <= 32'hFFFFFFFF;
                    11'h39A : DATO <= 32'hFFFFFFFF;
                    11'h39B : DATO <= 32'hFFFFFFFF;
                    11'h39C : DATO <= 32'hFFFFFFFF;
                    11'h39D : DATO <= 32'hFFFFFFFF;
                    11'h39E : DATO <= 32'hFFFFFFFF;
                    11'h39F : DATO <= 32'hFFFFFFFF;
                    11'h3A0 : DATO <= 32'hFFFFFFFF;
                    11'h3A1 : DATO <= 32'hFFFFFFFF;
                    11'h3A2 : DATO <= 32'hFFFFFFFF;
                    11'h3A3 : DATO <= 32'hFFFFFFFF;
                    11'h3A4 : DATO <= 32'hFFFFFFFF;
                    11'h3A5 : DATO <= 32'hFFFFFFFF;
                    11'h3A6 : DATO <= 32'hFFFFFFFF;
                    11'h3A7 : DATO <= 32'hFFFFFFFF;
                    11'h3A8 : DATO <= 32'hFFFFFFFF;
                    11'h3A9 : DATO <= 32'hFFFFFFFF;
                    11'h3AA : DATO <= 32'hFFFFFFFF;
                    11'h3AB : DATO <= 32'hFFFFFFFF;
                    11'h3AC : DATO <= 32'hFFFFFFFF;
                    11'h3AD : DATO <= 32'hFFFFFFFF;
                    11'h3AE : DATO <= 32'hFFFFFFFF;
                    11'h3AF : DATO <= 32'hFFFFFFFF;
                    11'h3B0 : DATO <= 32'hFFFFFFFF;
                    11'h3B1 : DATO <= 32'hFFFFFFFF;
                    11'h3B2 : DATO <= 32'hFFFFFFFF;
                    11'h3B3 : DATO <= 32'hFFFFFFFF;
                    11'h3B4 : DATO <= 32'hFFFFFFFF;
                    11'h3B5 : DATO <= 32'hFFFFFFFF;
                    11'h3B6 : DATO <= 32'hFFFFFFFF;
                    11'h3B7 : DATO <= 32'hFFFFFFFF;
                    11'h3B8 : DATO <= 32'hFFFFFFFF;
                    11'h3B9 : DATO <= 32'hFFFFFFFF;
                    11'h3BA : DATO <= 32'hFFFFFFFF;
                    11'h3BB : DATO <= 32'hFFFFFFFF;
                    11'h3BC : DATO <= 32'hFFFFFFFF;
                    11'h3BD : DATO <= 32'hFFFFFFFF;
                    11'h3BE : DATO <= 32'hFFFFFFFF;
                    11'h3BF : DATO <= 32'hFFFFFFFF;
                    11'h3C0 : DATO <= 32'hFFFFFFFF;
                    11'h3C1 : DATO <= 32'hFFFFFFFF;
                    11'h3C2 : DATO <= 32'hFFFFFFFF;
                    11'h3C3 : DATO <= 32'hFFFFFFFF;
                    11'h3C4 : DATO <= 32'hFFFFFFFF;
                    11'h3C5 : DATO <= 32'hFFFFFFFF;
                    11'h3C6 : DATO <= 32'hFFFFFFFF;
                    11'h3C7 : DATO <= 32'hFFFFFFFF;
                    11'h3C8 : DATO <= 32'hFFFFFFFF;
                    11'h3C9 : DATO <= 32'hFFFFFFFF;
                    11'h3CA : DATO <= 32'hFFFFFFFF;
                    11'h3CB : DATO <= 32'hFFFFFFFF;
                    11'h3CC : DATO <= 32'hFFFFFFFF;
                    11'h3CD : DATO <= 32'hFFFFFFFF;
                    11'h3CE : DATO <= 32'hFFFFFFFF;
                    11'h3CF : DATO <= 32'hFFFFFFFF;
                    11'h3D0 : DATO <= 32'hFFFFFFFF;
                    11'h3D1 : DATO <= 32'hFFFFFFFF;
                    11'h3D2 : DATO <= 32'hFFFFFFFF;
                    11'h3D3 : DATO <= 32'hFFFFFFFF;
                    11'h3D4 : DATO <= 32'hFFFFFFFF;
                    11'h3D5 : DATO <= 32'hFFFFFFFF;
                    11'h3D6 : DATO <= 32'hFFFFFFFF;
                    11'h3D7 : DATO <= 32'hFFFFFFFF;
                    11'h3D8 : DATO <= 32'hFFFFFFFF;
                    11'h3D9 : DATO <= 32'hFFFFFFFF;
                    11'h3DA : DATO <= 32'hFFFFFFFF;
                    11'h3DB : DATO <= 32'hFFFFFFFF;
                    11'h3DC : DATO <= 32'hFFFFFFFF;
                    11'h3DD : DATO <= 32'hFFFFFFFF;
                    11'h3DE : DATO <= 32'hFFFFFFFF;
                    11'h3DF : DATO <= 32'hFFFFFFFF;
                    11'h3E0 : DATO <= 32'hFFFFFFFF;
                    11'h3E1 : DATO <= 32'hFFFFFFFF;
                    11'h3E2 : DATO <= 32'hFFFFFFFF;
                    11'h3E3 : DATO <= 32'hFFFFFFFF;
                    11'h3E4 : DATO <= 32'hFFFFFFFF;
                    11'h3E5 : DATO <= 32'hFFFFFFFF;
                    11'h3E6 : DATO <= 32'hFFFFFFFF;
                    11'h3E7 : DATO <= 32'hFFFFFFFF;
                    11'h3E8 : DATO <= 32'hFFFFFFFF;
                    11'h3E9 : DATO <= 32'hFFFFFFFF;
                    11'h3EA : DATO <= 32'hFFFFFFFF;
                    11'h3EB : DATO <= 32'hFFFFFFFF;
                    11'h3EC : DATO <= 32'hFFFFFFFF;
                    11'h3ED : DATO <= 32'hFFFFFFFF;
                    11'h3EE : DATO <= 32'hFFFFFFFF;
                    11'h3EF : DATO <= 32'hFFFFFFFF;
                    11'h3F0 : DATO <= 32'hFFFFFFFF;
                    11'h3F1 : DATO <= 32'hFFFFFFFF;
                    11'h3F2 : DATO <= 32'hFFFFFFFF;
                    11'h3F3 : DATO <= 32'hFFFFFFFF;
                    11'h3F4 : DATO <= 32'hFFFFFFFF;
                    11'h3F5 : DATO <= 32'hFFFFFFFF;
                    11'h3F6 : DATO <= 32'hFFFFFFFF;
                    11'h3F7 : DATO <= 32'hFFFFFFFF;
                    11'h3F8 : DATO <= 32'hFFFFFFFF;
                    11'h3F9 : DATO <= 32'hFFFFFFFF;
                    11'h3FA : DATO <= 32'hFFFFFFFF;
                    11'h3FB : DATO <= 32'hFFFFFFFF;
                    11'h3FC : DATO <= 32'hFFFFFFFF;
                    11'h3FD : DATO <= 32'hFFFFFFFF;
                    11'h3FE : DATO <= 32'hFFFFFFFF;
                    11'h3FF : DATO <= 32'hFFFFFFFF;
                    11'h400 : DATO <= 32'hFFFFFFFF;
                    11'h401 : DATO <= 32'hFFFFFFFF;
                    11'h402 : DATO <= 32'hFFFFFFFF;
                    11'h403 : DATO <= 32'hFFFFFFFF;
                    11'h404 : DATO <= 32'hFFFFFFFF;
                    11'h405 : DATO <= 32'hFFFFFFFF;
                    11'h406 : DATO <= 32'hFFFFFFFF;
                    11'h407 : DATO <= 32'hFFFFFFFF;
                    11'h408 : DATO <= 32'hFFFFFFFF;
                    11'h409 : DATO <= 32'hFFFFFFFF;
                    11'h40A : DATO <= 32'hFFFFFFFF;
                    11'h40B : DATO <= 32'hFFFFFFFF;
                    11'h40C : DATO <= 32'hFFFFFFFF;
                    11'h40D : DATO <= 32'hFFFFFFFF;
                    11'h40E : DATO <= 32'hFFFFFFFF;
                    11'h40F : DATO <= 32'hFFFFFFFF;
                    11'h410 : DATO <= 32'hFFFFFFFF;
                    11'h411 : DATO <= 32'hFFFFFFFF;
                    11'h412 : DATO <= 32'hFFFFFFFF;
                    11'h413 : DATO <= 32'hFFFFFFFF;
                    11'h414 : DATO <= 32'hFFFFFFFF;
                    11'h415 : DATO <= 32'hFFFFFFFF;
                    11'h416 : DATO <= 32'hFFFFFFFF;
                    11'h417 : DATO <= 32'hFFFFFFFF;
                    11'h418 : DATO <= 32'hFFFFFFFF;
                    11'h419 : DATO <= 32'hFFFFFFFF;
                    11'h41A : DATO <= 32'hFFFFFFFF;
                    11'h41B : DATO <= 32'hFFFFFFFF;
                    11'h41C : DATO <= 32'hFFFFFFFF;
                    11'h41D : DATO <= 32'hFFFFFFFF;
                    11'h41E : DATO <= 32'hFFFFFFFF;
                    11'h41F : DATO <= 32'hFFFFFFFF;
                    11'h420 : DATO <= 32'hFFFFFFFF;
                    11'h421 : DATO <= 32'hFFFFFFFF;
                    11'h422 : DATO <= 32'hFFFFFFFF;
                    11'h423 : DATO <= 32'hFFFFFFFF;
                    11'h424 : DATO <= 32'hFFFFFFFF;
                    11'h425 : DATO <= 32'hFFFFFFFF;
                    11'h426 : DATO <= 32'hFFFFFFFF;
                    11'h427 : DATO <= 32'hFFFFFFFF;
                    11'h428 : DATO <= 32'hFFFFFFFF;
                    11'h429 : DATO <= 32'hFFFFFFFF;
                    11'h42A : DATO <= 32'hFFFFFFFF;
                    11'h42B : DATO <= 32'hFFFFFFFF;
                    11'h42C : DATO <= 32'hFFFFFFFF;
                    11'h42D : DATO <= 32'hFFFFFFFF;
                    11'h42E : DATO <= 32'hFFFFFFFF;
                    11'h42F : DATO <= 32'hFFFFFFFF;
                    11'h430 : DATO <= 32'hFFFFFFFF;
                    11'h431 : DATO <= 32'hFFFFFFFF;
                    11'h432 : DATO <= 32'hFFFFFFFF;
                    11'h433 : DATO <= 32'hFFFFFFFF;
                    11'h434 : DATO <= 32'hFFFFFFFF;
                    11'h435 : DATO <= 32'hFFFFFFFF;
                    11'h436 : DATO <= 32'hFFFFFFFF;
                    11'h437 : DATO <= 32'hFFFFFFFF;
                    11'h438 : DATO <= 32'hFFFFFFFF;
                    11'h439 : DATO <= 32'hFFFFFFFF;
                    11'h43A : DATO <= 32'hFFFFFFFF;
                    11'h43B : DATO <= 32'hFFFFFFFF;
                    11'h43C : DATO <= 32'hFFFFFFFF;
                    11'h43D : DATO <= 32'hFFFFFFFF;
                    11'h43E : DATO <= 32'hFFFFFFFF;
                    11'h43F : DATO <= 32'hFFFFFFFF;
                    11'h440 : DATO <= 32'hFFFFFFFF;
                    11'h441 : DATO <= 32'hFFFFFFFF;
                    11'h442 : DATO <= 32'hFFFFFFFF;
                    11'h443 : DATO <= 32'hFFFFFFFF;
                    11'h444 : DATO <= 32'hFFFFFFFF;
                    11'h445 : DATO <= 32'hFFFFFFFF;
                    11'h446 : DATO <= 32'hFFFFFFFF;
                    11'h447 : DATO <= 32'hFFFFFFFF;
                    11'h448 : DATO <= 32'hFFFFFFFF;
                    11'h449 : DATO <= 32'hFFFFFFFF;
                    11'h44A : DATO <= 32'hFFFFFFFF;
                    11'h44B : DATO <= 32'hFFFFFFFF;
                    11'h44C : DATO <= 32'hFFFFFFFF;
                    11'h44D : DATO <= 32'hFFFFFFFF;
                    11'h44E : DATO <= 32'hFFFFFFFF;
                    11'h44F : DATO <= 32'hFFFFFFFF;
                    11'h450 : DATO <= 32'hFFFFFFFF;
                    11'h451 : DATO <= 32'hFFFFFFFF;
                    11'h452 : DATO <= 32'hFFFFFFFF;
                    11'h453 : DATO <= 32'hFFFFFFFF;
                    11'h454 : DATO <= 32'hFFFFFFFF;
                    11'h455 : DATO <= 32'hFFFFFFFF;
                    11'h456 : DATO <= 32'hFFFFFFFF;
                    11'h457 : DATO <= 32'hFFFFFFFF;
                    11'h458 : DATO <= 32'hFFFFFFFF;
                    11'h459 : DATO <= 32'hFFFFFFFF;
                    11'h45A : DATO <= 32'hFFFFFFFF;
                    11'h45B : DATO <= 32'hFFFFFFFF;
                    11'h45C : DATO <= 32'hFFFFFFFF;
                    11'h45D : DATO <= 32'hFFFFFFFF;
                    11'h45E : DATO <= 32'hFFFFFFFF;
                    11'h45F : DATO <= 32'hFFFFFFFF;
                    11'h460 : DATO <= 32'hFFFFFFFF;
                    11'h461 : DATO <= 32'hFFFFFFFF;
                    11'h462 : DATO <= 32'hFFFFFFFF;
                    11'h463 : DATO <= 32'hFFFFFFFF;
                    11'h464 : DATO <= 32'hFFFFFFFF;
                    11'h465 : DATO <= 32'hFFFFFFFF;
                    11'h466 : DATO <= 32'hFFFFFFFF;
                    11'h467 : DATO <= 32'hFFFFFFFF;
                    11'h468 : DATO <= 32'hFFFFFFFF;
                    11'h469 : DATO <= 32'hFFFFFFFF;
                    11'h46A : DATO <= 32'hFFFFFFFF;
                    11'h46B : DATO <= 32'hFFFFFFFF;
                    11'h46C : DATO <= 32'hFFFFFFFF;
                    11'h46D : DATO <= 32'hFFFFFFFF;
                    11'h46E : DATO <= 32'hFFFFFFFF;
                    11'h46F : DATO <= 32'hFFFFFFFF;
                    11'h470 : DATO <= 32'hFFFFFFFF;
                    11'h471 : DATO <= 32'hFFFFFFFF;
                    11'h472 : DATO <= 32'hFFFFFFFF;
                    11'h473 : DATO <= 32'hFFFFFFFF;
                    11'h474 : DATO <= 32'hFFFFFFFF;
                    11'h475 : DATO <= 32'hFFFFFFFF;
                    11'h476 : DATO <= 32'hFFFFFFFF;
                    11'h477 : DATO <= 32'hFFFFFFFF;
                    11'h478 : DATO <= 32'hFFFFFFFF;
                    11'h479 : DATO <= 32'hFFFFFFFF;
                    11'h47A : DATO <= 32'hFFFFFFFF;
                    11'h47B : DATO <= 32'hFFFFFFFF;
                    11'h47C : DATO <= 32'hFFFFFFFF;
                    11'h47D : DATO <= 32'hFFFFFFFF;
                    11'h47E : DATO <= 32'hFFFFFFFF;
                    11'h47F : DATO <= 32'hFFFFFFFF;
                    11'h480 : DATO <= 32'hFFFFFFFF;
                    11'h481 : DATO <= 32'hFFFFFFFF;
                    11'h482 : DATO <= 32'hFFFFFFFF;
                    11'h483 : DATO <= 32'hFFFFFFFF;
                    11'h484 : DATO <= 32'hFFFFFFFF;
                    11'h485 : DATO <= 32'hFFFFFFFF;
                    11'h486 : DATO <= 32'hFFFFFFFF;
                    11'h487 : DATO <= 32'hFFFFFFFF;
                    11'h488 : DATO <= 32'hFFFFFFFF;
                    11'h489 : DATO <= 32'hFFFFFFFF;
                    11'h48A : DATO <= 32'hFFFFFFFF;
                    11'h48B : DATO <= 32'hFFFFFFFF;
                    11'h48C : DATO <= 32'hFFFFFFFF;
                    11'h48D : DATO <= 32'hFFFFFFFF;
                    11'h48E : DATO <= 32'hFFFFFFFF;
                    11'h48F : DATO <= 32'hFFFFFFFF;
                    11'h490 : DATO <= 32'hFFFFFFFF;
                    11'h491 : DATO <= 32'hFFFFFFFF;
                    11'h492 : DATO <= 32'hFFFFFFFF;
                    11'h493 : DATO <= 32'hFFFFFFFF;
                    11'h494 : DATO <= 32'hFFFFFFFF;
                    11'h495 : DATO <= 32'hFFFFFFFF;
                    11'h496 : DATO <= 32'hFFFFFFFF;
                    11'h497 : DATO <= 32'hFFFFFFFF;
                    11'h498 : DATO <= 32'hFFFFFFFF;
                    11'h499 : DATO <= 32'hFFFFFFFF;
                    11'h49A : DATO <= 32'hFFFFFFFF;
                    11'h49B : DATO <= 32'hFFFFFFFF;
                    11'h49C : DATO <= 32'hFFFFFFFF;
                    11'h49D : DATO <= 32'hFFFFFFFF;
                    11'h49E : DATO <= 32'hFFFFFFFF;
                    11'h49F : DATO <= 32'hFFFFFFFF;
                    11'h4A0 : DATO <= 32'hFFFFFFFF;
                    11'h4A1 : DATO <= 32'hFFFFFFFF;
                    11'h4A2 : DATO <= 32'hFFFFFFFF;
                    11'h4A3 : DATO <= 32'hFFFFFFFF;
                    11'h4A4 : DATO <= 32'hFFFFFFFF;
                    11'h4A5 : DATO <= 32'hFFFFFFFF;
                    11'h4A6 : DATO <= 32'hFFFFFFFF;
                    11'h4A7 : DATO <= 32'hFFFFFFFF;
                    11'h4A8 : DATO <= 32'hFFFFFFFF;
                    11'h4A9 : DATO <= 32'hFFFFFFFF;
                    11'h4AA : DATO <= 32'hFFFFFFFF;
                    11'h4AB : DATO <= 32'hFFFFFFFF;
                    11'h4AC : DATO <= 32'hFFFFFFFF;
                    11'h4AD : DATO <= 32'hFFFFFFFF;
                    11'h4AE : DATO <= 32'hFFFFFFFF;
                    11'h4AF : DATO <= 32'hFFFFFFFF;
                    11'h4B0 : DATO <= 32'hFFFFFFFF;
                    11'h4B1 : DATO <= 32'hFFFFFFFF;
                    11'h4B2 : DATO <= 32'hFFFFFFFF;
                    11'h4B3 : DATO <= 32'hFFFFFFFF;
                    11'h4B4 : DATO <= 32'hFFFFFFFF;
                    11'h4B5 : DATO <= 32'hFFFFFFFF;
                    11'h4B6 : DATO <= 32'hFFFFFFFF;
                    11'h4B7 : DATO <= 32'hFFFFFFFF;
                    11'h4B8 : DATO <= 32'hFFFFFFFF;
                    11'h4B9 : DATO <= 32'hFFFFFFFF;
                    11'h4BA : DATO <= 32'hFFFFFFFF;
                    11'h4BB : DATO <= 32'hFFFFFFFF;
                    11'h4BC : DATO <= 32'hFFFFFFFF;
                    11'h4BD : DATO <= 32'hFFFFFFFF;
                    11'h4BE : DATO <= 32'hFFFFFFFF;
                    11'h4BF : DATO <= 32'hFFFFFFFF;
                    11'h4C0 : DATO <= 32'hFFFFFFFF;
                    11'h4C1 : DATO <= 32'hFFFFFFFF;
                    11'h4C2 : DATO <= 32'hFFFFFFFF;
                    11'h4C3 : DATO <= 32'hFFFFFFFF;
                    11'h4C4 : DATO <= 32'hFFFFFFFF;
                    11'h4C5 : DATO <= 32'hFFFFFFFF;
                    11'h4C6 : DATO <= 32'hFFFFFFFF;
                    11'h4C7 : DATO <= 32'hFFFFFFFF;
                    11'h4C8 : DATO <= 32'hFFFFFFFF;
                    11'h4C9 : DATO <= 32'hFFFFFFFF;
                    11'h4CA : DATO <= 32'hFFFFFFFF;
                    11'h4CB : DATO <= 32'hFFFFFFFF;
                    11'h4CC : DATO <= 32'hFFFFFFFF;
                    11'h4CD : DATO <= 32'hFFFFFFFF;
                    11'h4CE : DATO <= 32'hFFFFFFFF;
                    11'h4CF : DATO <= 32'hFFFFFFFF;
                    11'h4D0 : DATO <= 32'hFFFFFFFF;
                    11'h4D1 : DATO <= 32'hFFFFFFFF;
                    11'h4D2 : DATO <= 32'hFFFFFFFF;
                    11'h4D3 : DATO <= 32'hFFFFFFFF;
                    11'h4D4 : DATO <= 32'hFFFFFFFF;
                    11'h4D5 : DATO <= 32'hFFFFFFFF;
                    11'h4D6 : DATO <= 32'hFFFFFFFF;
                    11'h4D7 : DATO <= 32'hFFFFFFFF;
                    11'h4D8 : DATO <= 32'hFFFFFFFF;
                    11'h4D9 : DATO <= 32'hFFFFFFFF;
                    11'h4DA : DATO <= 32'hFFFFFFFF;
                    11'h4DB : DATO <= 32'hFFFFFFFF;
                    11'h4DC : DATO <= 32'hFFFFFFFF;
                    11'h4DD : DATO <= 32'hFFFFFFFF;
                    11'h4DE : DATO <= 32'hFFFFFFFF;
                    11'h4DF : DATO <= 32'hFFFFFFFF;
                    11'h4E0 : DATO <= 32'hFFFFFFFF;
                    11'h4E1 : DATO <= 32'hFFFFFFFF;
                    11'h4E2 : DATO <= 32'hFFFFFFFF;
                    11'h4E3 : DATO <= 32'hFFFFFFFF;
                    11'h4E4 : DATO <= 32'hFFFFFFFF;
                    11'h4E5 : DATO <= 32'hFFFFFFFF;
                    11'h4E6 : DATO <= 32'hFFFFFFFF;
                    11'h4E7 : DATO <= 32'hFFFFFFFF;
                    11'h4E8 : DATO <= 32'hFFFFFFFF;
                    11'h4E9 : DATO <= 32'hFFFFFFFF;
                    11'h4EA : DATO <= 32'hFFFFFFFF;
                    11'h4EB : DATO <= 32'hFFFFFFFF;
                    11'h4EC : DATO <= 32'hFFFFFFFF;
                    11'h4ED : DATO <= 32'hFFFFFFFF;
                    11'h4EE : DATO <= 32'hFFFFFFFF;
                    11'h4EF : DATO <= 32'hFFFFFFFF;
                    11'h4F0 : DATO <= 32'hFFFFFFFF;
                    11'h4F1 : DATO <= 32'hFFFFFFFF;
                    11'h4F2 : DATO <= 32'hFFFFFFFF;
                    11'h4F3 : DATO <= 32'hFFFFFFFF;
                    11'h4F4 : DATO <= 32'hFFFFFFFF;
                    11'h4F5 : DATO <= 32'hFFFFFFFF;
                    11'h4F6 : DATO <= 32'hFFFFFFFF;
                    11'h4F7 : DATO <= 32'hFFFFFFFF;
                    11'h4F8 : DATO <= 32'hFFFFFFFF;
                    11'h4F9 : DATO <= 32'hFFFFFFFF;
                    11'h4FA : DATO <= 32'hFFFFFFFF;
                    11'h4FB : DATO <= 32'hFFFFFFFF;
                    11'h4FC : DATO <= 32'hFFFFFFFF;
                    11'h4FD : DATO <= 32'hFFFFFFFF;
                    11'h4FE : DATO <= 32'hFFFFFFFF;
                    11'h4FF : DATO <= 32'hFFFFFFFF;
                    11'h500 : DATO <= 32'hFFFFFFFF;
                    11'h501 : DATO <= 32'hFFFFFFFF;
                    11'h502 : DATO <= 32'hFFFFFFFF;
                    11'h503 : DATO <= 32'hFFFFFFFF;
                    11'h504 : DATO <= 32'hFFFFFFFF;
                    11'h505 : DATO <= 32'hFFFFFFFF;
                    11'h506 : DATO <= 32'hFFFFFFFF;
                    11'h507 : DATO <= 32'hFFFFFFFF;
                    11'h508 : DATO <= 32'hFFFFFFFF;
                    11'h509 : DATO <= 32'hFFFFFFFF;
                    11'h50A : DATO <= 32'hFFFFFFFF;
                    11'h50B : DATO <= 32'hFFFFFFFF;
                    11'h50C : DATO <= 32'hFFFFFFFF;
                    11'h50D : DATO <= 32'hFFFFFFFF;
                    11'h50E : DATO <= 32'hFFFFFFFF;
                    11'h50F : DATO <= 32'hFFFFFFFF;
                    11'h510 : DATO <= 32'hFFFFFFFF;
                    11'h511 : DATO <= 32'hFFFFFFFF;
                    11'h512 : DATO <= 32'hFFFFFFFF;
                    11'h513 : DATO <= 32'hFFFFFFFF;
                    11'h514 : DATO <= 32'hFFFFFFFF;
                    11'h515 : DATO <= 32'hFFFFFFFF;
                    11'h516 : DATO <= 32'hFFFFFFFF;
                    11'h517 : DATO <= 32'hFFFFFFFF;
                    11'h518 : DATO <= 32'hFFFFFFFF;
                    11'h519 : DATO <= 32'hFFFFFFFF;
                    11'h51A : DATO <= 32'hFFFFFFFF;
                    11'h51B : DATO <= 32'hFFFFFFFF;
                    11'h51C : DATO <= 32'hFFFFFFFF;
                    11'h51D : DATO <= 32'hFFFFFFFF;
                    11'h51E : DATO <= 32'hFFFFFFFF;
                    11'h51F : DATO <= 32'hFFFFFFFF;
                    11'h520 : DATO <= 32'hFFFFFFFF;
                    11'h521 : DATO <= 32'hFFFFFFFF;
                    11'h522 : DATO <= 32'hFFFFFFFF;
                    11'h523 : DATO <= 32'hFFFFFFFF;
                    11'h524 : DATO <= 32'hFFFFFFFF;
                    11'h525 : DATO <= 32'hFFFFFFFF;
                    11'h526 : DATO <= 32'hFFFFFFFF;
                    11'h527 : DATO <= 32'hFFFFFFFF;
                    11'h528 : DATO <= 32'hFFFFFFFF;
                    11'h529 : DATO <= 32'hFFFFFFFF;
                    11'h52A : DATO <= 32'hFFFFFFFF;
                    11'h52B : DATO <= 32'hFFFFFFFF;
                    11'h52C : DATO <= 32'hFFFFFFFF;
                    11'h52D : DATO <= 32'hFFFFFFFF;
                    11'h52E : DATO <= 32'hFFFFFFFF;
                    11'h52F : DATO <= 32'hFFFFFFFF;
                    11'h530 : DATO <= 32'hFFFFFFFF;
                    11'h531 : DATO <= 32'hFFFFFFFF;
                    11'h532 : DATO <= 32'hFFFFFFFF;
                    11'h533 : DATO <= 32'hFFFFFFFF;
                    11'h534 : DATO <= 32'hFFFFFFFF;
                    11'h535 : DATO <= 32'hFFFFFFFF;
                    11'h536 : DATO <= 32'hFFFFFFFF;
                    11'h537 : DATO <= 32'hFFFFFFFF;
                    11'h538 : DATO <= 32'hFFFFFFFF;
                    11'h539 : DATO <= 32'hFFFFFFFF;
                    11'h53A : DATO <= 32'hFFFFFFFF;
                    11'h53B : DATO <= 32'hFFFFFFFF;
                    11'h53C : DATO <= 32'hFFFFFFFF;
                    11'h53D : DATO <= 32'hFFFFFFFF;
                    11'h53E : DATO <= 32'hFFFFFFFF;
                    11'h53F : DATO <= 32'hFFFFFFFF;
                    11'h540 : DATO <= 32'hFFFFFFFF;
                    11'h541 : DATO <= 32'hFFFFFFFF;
                    11'h542 : DATO <= 32'hFFFFFFFF;
                    11'h543 : DATO <= 32'hFFFFFFFF;
                    11'h544 : DATO <= 32'hFFFFFFFF;
                    11'h545 : DATO <= 32'hFFFFFFFF;
                    11'h546 : DATO <= 32'hFFFFFFFF;
                    11'h547 : DATO <= 32'hFFFFFFFF;
                    11'h548 : DATO <= 32'hFFFFFFFF;
                    11'h549 : DATO <= 32'hFFFFFFFF;
                    11'h54A : DATO <= 32'hFFFFFFFF;
                    11'h54B : DATO <= 32'hFFFFFFFF;
                    11'h54C : DATO <= 32'hFFFFFFFF;
                    11'h54D : DATO <= 32'hFFFFFFFF;
                    11'h54E : DATO <= 32'hFFFFFFFF;
                    11'h54F : DATO <= 32'hFFFFFFFF;
                    11'h550 : DATO <= 32'hFFFFFFFF;
                    11'h551 : DATO <= 32'hFFFFFFFF;
                    11'h552 : DATO <= 32'hFFFFFFFF;
                    11'h553 : DATO <= 32'hFFFFFFFF;
                    11'h554 : DATO <= 32'hFFFFFFFF;
                    11'h555 : DATO <= 32'hFFFFFFFF;
                    11'h556 : DATO <= 32'hFFFFFFFF;
                    11'h557 : DATO <= 32'hFFFFFFFF;
                    11'h558 : DATO <= 32'hFFFFFFFF;
                    11'h559 : DATO <= 32'hFFFFFFFF;
                    11'h55A : DATO <= 32'hFFFFFFFF;
                    11'h55B : DATO <= 32'hFFFFFFFF;
                    11'h55C : DATO <= 32'hFFFFFFFF;
                    11'h55D : DATO <= 32'hFFFFFFFF;
                    11'h55E : DATO <= 32'hFFFFFFFF;
                    11'h55F : DATO <= 32'hFFFFFFFF;
                    11'h560 : DATO <= 32'hFFFFFFFF;
                    11'h561 : DATO <= 32'hFFFFFFFF;
                    11'h562 : DATO <= 32'hFFFFFFFF;
                    11'h563 : DATO <= 32'hFFFFFFFF;
                    11'h564 : DATO <= 32'hFFFFFFFF;
                    11'h565 : DATO <= 32'hFFFFFFFF;
                    11'h566 : DATO <= 32'hFFFFFFFF;
                    11'h567 : DATO <= 32'hFFFFFFFF;
                    11'h568 : DATO <= 32'hFFFFFFFF;
                    11'h569 : DATO <= 32'hFFFFFFFF;
                    11'h56A : DATO <= 32'hFFFFFFFF;
                    11'h56B : DATO <= 32'hFFFFFFFF;
                    11'h56C : DATO <= 32'hFFFFFFFF;
                    11'h56D : DATO <= 32'hFFFFFFFF;
                    11'h56E : DATO <= 32'hFFFFFFFF;
                    11'h56F : DATO <= 32'hFFFFFFFF;
                    11'h570 : DATO <= 32'hFFFFFFFF;
                    11'h571 : DATO <= 32'hFFFFFFFF;
                    11'h572 : DATO <= 32'hFFFFFFFF;
                    11'h573 : DATO <= 32'hFFFFFFFF;
                    11'h574 : DATO <= 32'hFFFFFFFF;
                    11'h575 : DATO <= 32'hFFFFFFFF;
                    11'h576 : DATO <= 32'hFFFFFFFF;
                    11'h577 : DATO <= 32'hFFFFFFFF;
                    11'h578 : DATO <= 32'hFFFFFFFF;
                    11'h579 : DATO <= 32'hFFFFFFFF;
                    11'h57A : DATO <= 32'hFFFFFFFF;
                    11'h57B : DATO <= 32'hFFFFFFFF;
                    11'h57C : DATO <= 32'hFFFFFFFF;
                    11'h57D : DATO <= 32'hFFFFFFFF;
                    11'h57E : DATO <= 32'hFFFFFFFF;
                    11'h57F : DATO <= 32'hFFFFFFFF;
                    11'h580 : DATO <= 32'hFFFFFFFF;
                    11'h581 : DATO <= 32'hFFFFFFFF;
                    11'h582 : DATO <= 32'hFFFFFFFF;
                    11'h583 : DATO <= 32'hFFFFFFFF;
                    11'h584 : DATO <= 32'hFFFFFFFF;
                    11'h585 : DATO <= 32'hFFFFFFFF;
                    11'h586 : DATO <= 32'hFFFFFFFF;
                    11'h587 : DATO <= 32'hFFFFFFFF;
                    11'h588 : DATO <= 32'hFFFFFFFF;
                    11'h589 : DATO <= 32'hFFFFFFFF;
                    11'h58A : DATO <= 32'hFFFFFFFF;
                    11'h58B : DATO <= 32'hFFFFFFFF;
                    11'h58C : DATO <= 32'hFFFFFFFF;
                    11'h58D : DATO <= 32'hFFFFFFFF;
                    11'h58E : DATO <= 32'hFFFFFFFF;
                    11'h58F : DATO <= 32'hFFFFFFFF;
                    11'h590 : DATO <= 32'hFFFFFFFF;
                    11'h591 : DATO <= 32'hFFFFFFFF;
                    11'h592 : DATO <= 32'hFFFFFFFF;
                    11'h593 : DATO <= 32'hFFFFFFFF;
                    11'h594 : DATO <= 32'hFFFFFFFF;
                    11'h595 : DATO <= 32'hFFFFFFFF;
                    11'h596 : DATO <= 32'hFFFFFFFF;
                    11'h597 : DATO <= 32'hFFFFFFFF;
                    11'h598 : DATO <= 32'hFFFFFFFF;
                    11'h599 : DATO <= 32'hFFFFFFFF;
                    11'h59A : DATO <= 32'hFFFFFFFF;
                    11'h59B : DATO <= 32'hFFFFFFFF;
                    11'h59C : DATO <= 32'hFFFFFFFF;
                    11'h59D : DATO <= 32'hFFFFFFFF;
                    11'h59E : DATO <= 32'hFFFFFFFF;
                    11'h59F : DATO <= 32'hFFFFFFFF;
                    11'h5A0 : DATO <= 32'hFFFFFFFF;
                    11'h5A1 : DATO <= 32'hFFFFFFFF;
                    11'h5A2 : DATO <= 32'hFFFFFFFF;
                    11'h5A3 : DATO <= 32'hFFFFFFFF;
                    11'h5A4 : DATO <= 32'hFFFFFFFF;
                    11'h5A5 : DATO <= 32'hFFFFFFFF;
                    11'h5A6 : DATO <= 32'hFFFFFFFF;
                    11'h5A7 : DATO <= 32'hFFFFFFFF;
                    11'h5A8 : DATO <= 32'hFFFFFFFF;
                    11'h5A9 : DATO <= 32'hFFFFFFFF;
                    11'h5AA : DATO <= 32'hFFFFFFFF;
                    11'h5AB : DATO <= 32'hFFFFFFFF;
                    11'h5AC : DATO <= 32'hFFFFFFFF;
                    11'h5AD : DATO <= 32'hFFFFFFFF;
                    11'h5AE : DATO <= 32'hFFFFFFFF;
                    11'h5AF : DATO <= 32'hFFFFFFFF;
                    11'h5B0 : DATO <= 32'hFFFFFFFF;
                    11'h5B1 : DATO <= 32'hFFFFFFFF;
                    11'h5B2 : DATO <= 32'hFFFFFFFF;
                    11'h5B3 : DATO <= 32'hFFFFFFFF;
                    11'h5B4 : DATO <= 32'hFFFFFFFF;
                    11'h5B5 : DATO <= 32'hFFFFFFFF;
                    11'h5B6 : DATO <= 32'hFFFFFFFF;
                    11'h5B7 : DATO <= 32'hFFFFFFFF;
                    11'h5B8 : DATO <= 32'hFFFFFFFF;
                    11'h5B9 : DATO <= 32'hFFFFFFFF;
                    11'h5BA : DATO <= 32'hFFFFFFFF;
                    11'h5BB : DATO <= 32'hFFFFFFFF;
                    11'h5BC : DATO <= 32'hFFFFFFFF;
                    11'h5BD : DATO <= 32'hFFFFFFFF;
                    11'h5BE : DATO <= 32'hFFFFFFFF;
                    11'h5BF : DATO <= 32'hFFFFFFFF;
                    11'h5C0 : DATO <= 32'hFFFFFFFF;
                    11'h5C1 : DATO <= 32'hFFFFFFFF;
                    11'h5C2 : DATO <= 32'hFFFFFFFF;
                    11'h5C3 : DATO <= 32'hFFFFFFFF;
                    11'h5C4 : DATO <= 32'hFFFFFFFF;
                    11'h5C5 : DATO <= 32'hFFFFFFFF;
                    11'h5C6 : DATO <= 32'hFFFFFFFF;
                    11'h5C7 : DATO <= 32'hFFFFFFFF;
                    11'h5C8 : DATO <= 32'hFFFFFFFF;
                    11'h5C9 : DATO <= 32'hFFFFFFFF;
                    11'h5CA : DATO <= 32'hFFFFFFFF;
                    11'h5CB : DATO <= 32'hFFFFFFFF;
                    11'h5CC : DATO <= 32'hFFFFFFFF;
                    11'h5CD : DATO <= 32'hFFFFFFFF;
                    11'h5CE : DATO <= 32'hFFFFFFFF;
                    11'h5CF : DATO <= 32'hFFFFFFFF;
                    11'h5D0 : DATO <= 32'hFFFFFFFF;
                    11'h5D1 : DATO <= 32'hFFFFFFFF;
                    11'h5D2 : DATO <= 32'hFFFFFFFF;
                    11'h5D3 : DATO <= 32'hFFFFFFFF;
                    11'h5D4 : DATO <= 32'hFFFFFFFF;
                    11'h5D5 : DATO <= 32'hFFFFFFFF;
                    11'h5D6 : DATO <= 32'hFFFFFFFF;
                    11'h5D7 : DATO <= 32'hFFFFFFFF;
                    11'h5D8 : DATO <= 32'hFFFFFFFF;
                    11'h5D9 : DATO <= 32'hFFFFFFFF;
                    11'h5DA : DATO <= 32'hFFFFFFFF;
                    11'h5DB : DATO <= 32'hFFFFFFFF;
                    11'h5DC : DATO <= 32'hFFFFFFFF;
                    11'h5DD : DATO <= 32'hFFFFFFFF;
                    11'h5DE : DATO <= 32'hFFFFFFFF;
                    11'h5DF : DATO <= 32'hFFFFFFFF;
                    11'h5E0 : DATO <= 32'hFFFFFFFF;
                    11'h5E1 : DATO <= 32'hFFFFFFFF;
                    11'h5E2 : DATO <= 32'hFFFFFFFF;
                    11'h5E3 : DATO <= 32'hFFFFFFFF;
                    11'h5E4 : DATO <= 32'hFFFFFFFF;
                    11'h5E5 : DATO <= 32'hFFFFFFFF;
                    11'h5E6 : DATO <= 32'hFFFFFFFF;
                    11'h5E7 : DATO <= 32'hFFFFFFFF;
                    11'h5E8 : DATO <= 32'hFFFFFFFF;
                    11'h5E9 : DATO <= 32'hFFFFFFFF;
                    11'h5EA : DATO <= 32'hFFFFFFFF;
                    11'h5EB : DATO <= 32'hFFFFFFFF;
                    11'h5EC : DATO <= 32'hFFFFFFFF;
                    11'h5ED : DATO <= 32'hFFFFFFFF;
                    11'h5EE : DATO <= 32'hFFFFFFFF;
                    11'h5EF : DATO <= 32'hFFFFFFFF;
                    11'h5F0 : DATO <= 32'hFFFFFFFF;
                    11'h5F1 : DATO <= 32'hFFFFFFFF;
                    11'h5F2 : DATO <= 32'hFFFFFFFF;
                    11'h5F3 : DATO <= 32'hFFFFFFFF;
                    11'h5F4 : DATO <= 32'hFFFFFFFF;
                    11'h5F5 : DATO <= 32'hFFFFFFFF;
                    11'h5F6 : DATO <= 32'hFFFFFFFF;
                    11'h5F7 : DATO <= 32'hFFFFFFFF;
                    11'h5F8 : DATO <= 32'hFFFFFFFF;
                    11'h5F9 : DATO <= 32'hFFFFFFFF;
                    11'h5FA : DATO <= 32'hFFFFFFFF;
                    11'h5FB : DATO <= 32'hFFFFFFFF;
                    11'h5FC : DATO <= 32'hFFFFFFFF;
                    11'h5FD : DATO <= 32'hFFFFFFFF;
                    11'h5FE : DATO <= 32'hFFFFFFFF;
                    11'h5FF : DATO <= 32'hFFFFFFFF;
                    11'h600 : DATO <= 32'hFFFFFFFF;
                    11'h601 : DATO <= 32'hFFFFFFFF;
                    11'h602 : DATO <= 32'hFFFFFFFF;
                    11'h603 : DATO <= 32'hFFFFFFFF;
                    11'h604 : DATO <= 32'hFFFFFFFF;
                    11'h605 : DATO <= 32'hFFFFFFFF;
                    11'h606 : DATO <= 32'hFFFFFFFF;
                    11'h607 : DATO <= 32'hFFFFFFFF;
                    11'h608 : DATO <= 32'hFFFFFFFF;
                    11'h609 : DATO <= 32'hFFFFFFFF;
                    11'h60A : DATO <= 32'hFFFFFFFF;
                    11'h60B : DATO <= 32'hFFFFFFFF;
                    11'h60C : DATO <= 32'hFFFFFFFF;
                    11'h60D : DATO <= 32'hFFFFFFFF;
                    11'h60E : DATO <= 32'hFFFFFFFF;
                    11'h60F : DATO <= 32'hFFFFFFFF;
                    11'h610 : DATO <= 32'hFFFFFFFF;
                    11'h611 : DATO <= 32'hFFFFFFFF;
                    11'h612 : DATO <= 32'hFFFFFFFF;
                    11'h613 : DATO <= 32'hFFFFFFFF;
                    11'h614 : DATO <= 32'hFFFFFFFF;
                    11'h615 : DATO <= 32'hFFFFFFFF;
                    11'h616 : DATO <= 32'hFFFFFFFF;
                    11'h617 : DATO <= 32'hFFFFFFFF;
                    11'h618 : DATO <= 32'hFFFFFFFF;
                    11'h619 : DATO <= 32'hFFFFFFFF;
                    11'h61A : DATO <= 32'hFFFFFFFF;
                    11'h61B : DATO <= 32'hFFFFFFFF;
                    11'h61C : DATO <= 32'hFFFFFFFF;
                    11'h61D : DATO <= 32'hFFFFFFFF;
                    11'h61E : DATO <= 32'hFFFFFFFF;
                    11'h61F : DATO <= 32'hFFFFFFFF;
                    11'h620 : DATO <= 32'hFFFFFFFF;
                    11'h621 : DATO <= 32'hFFFFFFFF;
                    11'h622 : DATO <= 32'hFFFFFFFF;
                    11'h623 : DATO <= 32'hFFFFFFFF;
                    11'h624 : DATO <= 32'hFFFFFFFF;
                    11'h625 : DATO <= 32'hFFFFFFFF;
                    11'h626 : DATO <= 32'hFFFFFFFF;
                    11'h627 : DATO <= 32'hFFFFFFFF;
                    11'h628 : DATO <= 32'hFFFFFFFF;
                    11'h629 : DATO <= 32'hFFFFFFFF;
                    11'h62A : DATO <= 32'hFFFFFFFF;
                    11'h62B : DATO <= 32'hFFFFFFFF;
                    11'h62C : DATO <= 32'hFFFFFFFF;
                    11'h62D : DATO <= 32'hFFFFFFFF;
                    11'h62E : DATO <= 32'hFFFFFFFF;
                    11'h62F : DATO <= 32'hFFFFFFFF;
                    11'h630 : DATO <= 32'hFFFFFFFF;
                    11'h631 : DATO <= 32'hFFFFFFFF;
                    11'h632 : DATO <= 32'hFFFFFFFF;
                    11'h633 : DATO <= 32'hFFFFFFFF;
                    11'h634 : DATO <= 32'hFFFFFFFF;
                    11'h635 : DATO <= 32'hFFFFFFFF;
                    11'h636 : DATO <= 32'hFFFFFFFF;
                    11'h637 : DATO <= 32'hFFFFFFFF;
                    11'h638 : DATO <= 32'hFFFFFFFF;
                    11'h639 : DATO <= 32'hFFFFFFFF;
                    11'h63A : DATO <= 32'hFFFFFFFF;
                    11'h63B : DATO <= 32'hFFFFFFFF;
                    11'h63C : DATO <= 32'hFFFFFFFF;
                    11'h63D : DATO <= 32'hFFFFFFFF;
                    11'h63E : DATO <= 32'hFFFFFFFF;
                    11'h63F : DATO <= 32'hFFFFFFFF;
                    11'h640 : DATO <= 32'hFFFFFFFF;
                    11'h641 : DATO <= 32'hFFFFFFFF;
                    11'h642 : DATO <= 32'hFFFFFFFF;
                    11'h643 : DATO <= 32'hFFFFFFFF;
                    11'h644 : DATO <= 32'hFFFFFFFF;
                    11'h645 : DATO <= 32'hFFFFFFFF;
                    11'h646 : DATO <= 32'hFFFFFFFF;
                    11'h647 : DATO <= 32'hFFFFFFFF;
                    11'h648 : DATO <= 32'hFFFFFFFF;
                    11'h649 : DATO <= 32'hFFFFFFFF;
                    11'h64A : DATO <= 32'hFFFFFFFF;
                    11'h64B : DATO <= 32'hFFFFFFFF;
                    11'h64C : DATO <= 32'hFFFFFFFF;
                    11'h64D : DATO <= 32'hFFFFFFFF;
                    11'h64E : DATO <= 32'hFFFFFFFF;
                    11'h64F : DATO <= 32'hFFFFFFFF;
                    11'h650 : DATO <= 32'hFFFFFFFF;
                    11'h651 : DATO <= 32'hFFFFFFFF;
                    11'h652 : DATO <= 32'hFFFFFFFF;
                    11'h653 : DATO <= 32'hFFFFFFFF;
                    11'h654 : DATO <= 32'hFFFFFFFF;
                    11'h655 : DATO <= 32'hFFFFFFFF;
                    11'h656 : DATO <= 32'hFFFFFFFF;
                    11'h657 : DATO <= 32'hFFFFFFFF;
                    11'h658 : DATO <= 32'hFFFFFFFF;
                    11'h659 : DATO <= 32'hFFFFFFFF;
                    11'h65A : DATO <= 32'hFFFFFFFF;
                    11'h65B : DATO <= 32'hFFFFFFFF;
                    11'h65C : DATO <= 32'hFFFFFFFF;
                    11'h65D : DATO <= 32'hFFFFFFFF;
                    11'h65E : DATO <= 32'hFFFFFFFF;
                    11'h65F : DATO <= 32'hFFFFFFFF;
                    11'h660 : DATO <= 32'hFFFFFFFF;
                    11'h661 : DATO <= 32'hFFFFFFFF;
                    11'h662 : DATO <= 32'hFFFFFFFF;
                    11'h663 : DATO <= 32'hFFFFFFFF;
                    11'h664 : DATO <= 32'hFFFFFFFF;
                    11'h665 : DATO <= 32'hFFFFFFFF;
                    11'h666 : DATO <= 32'hFFFFFFFF;
                    11'h667 : DATO <= 32'hFFFFFFFF;
                    11'h668 : DATO <= 32'hFFFFFFFF;
                    11'h669 : DATO <= 32'hFFFFFFFF;
                    11'h66A : DATO <= 32'hFFFFFFFF;
                    11'h66B : DATO <= 32'hFFFFFFFF;
                    11'h66C : DATO <= 32'hFFFFFFFF;
                    11'h66D : DATO <= 32'hFFFFFFFF;
                    11'h66E : DATO <= 32'hFFFFFFFF;
                    11'h66F : DATO <= 32'hFFFFFFFF;
                    11'h670 : DATO <= 32'hFFFFFFFF;
                    11'h671 : DATO <= 32'hFFFFFFFF;
                    11'h672 : DATO <= 32'hFFFFFFFF;
                    11'h673 : DATO <= 32'hFFFFFFFF;
                    11'h674 : DATO <= 32'hFFFFFFFF;
                    11'h675 : DATO <= 32'hFFFFFFFF;
                    11'h676 : DATO <= 32'hFFFFFFFF;
                    11'h677 : DATO <= 32'hFFFFFFFF;
                    11'h678 : DATO <= 32'hFFFFFFFF;
                    11'h679 : DATO <= 32'hFFFFFFFF;
                    11'h67A : DATO <= 32'hFFFFFFFF;
                    11'h67B : DATO <= 32'hFFFFFFFF;
                    11'h67C : DATO <= 32'hFFFFFFFF;
                    11'h67D : DATO <= 32'hFFFFFFFF;
                    11'h67E : DATO <= 32'hFFFFFFFF;
                    11'h67F : DATO <= 32'hFFFFFFFF;
                    11'h680 : DATO <= 32'hFFFFFFFF;
                    11'h681 : DATO <= 32'hFFFFFFFF;
                    11'h682 : DATO <= 32'hFFFFFFFF;
                    11'h683 : DATO <= 32'hFFFFFFFF;
                    11'h684 : DATO <= 32'hFFFFFFFF;
                    11'h685 : DATO <= 32'hFFFFFFFF;
                    11'h686 : DATO <= 32'hFFFFFFFF;
                    11'h687 : DATO <= 32'hFFFFFFFF;
                    11'h688 : DATO <= 32'hFFFFFFFF;
                    11'h689 : DATO <= 32'hFFFFFFFF;
                    11'h68A : DATO <= 32'hFFFFFFFF;
                    11'h68B : DATO <= 32'hFFFFFFFF;
                    11'h68C : DATO <= 32'hFFFFFFFF;
                    11'h68D : DATO <= 32'hFFFFFFFF;
                    11'h68E : DATO <= 32'hFFFFFFFF;
                    11'h68F : DATO <= 32'hFFFFFFFF;
                    11'h690 : DATO <= 32'hFFFFFFFF;
                    11'h691 : DATO <= 32'hFFFFFFFF;
                    11'h692 : DATO <= 32'hFFFFFFFF;
                    11'h693 : DATO <= 32'hFFFFFFFF;
                    11'h694 : DATO <= 32'hFFFFFFFF;
                    11'h695 : DATO <= 32'hFFFFFFFF;
                    11'h696 : DATO <= 32'hFFFFFFFF;
                    11'h697 : DATO <= 32'hFFFFFFFF;
                    11'h698 : DATO <= 32'hFFFFFFFF;
                    11'h699 : DATO <= 32'hFFFFFFFF;
                    11'h69A : DATO <= 32'hFFFFFFFF;
                    11'h69B : DATO <= 32'hFFFFFFFF;
                    11'h69C : DATO <= 32'hFFFFFFFF;
                    11'h69D : DATO <= 32'hFFFFFFFF;
                    11'h69E : DATO <= 32'hFFFFFFFF;
                    11'h69F : DATO <= 32'hFFFFFFFF;
                    11'h6A0 : DATO <= 32'hFFFFFFFF;
                    11'h6A1 : DATO <= 32'hFFFFFFFF;
                    11'h6A2 : DATO <= 32'hFFFFFFFF;
                    11'h6A3 : DATO <= 32'hFFFFFFFF;
                    11'h6A4 : DATO <= 32'hFFFFFFFF;
                    11'h6A5 : DATO <= 32'hFFFFFFFF;
                    11'h6A6 : DATO <= 32'hFFFFFFFF;
                    11'h6A7 : DATO <= 32'hFFFFFFFF;
                    11'h6A8 : DATO <= 32'hFFFFFFFF;
                    11'h6A9 : DATO <= 32'hFFFFFFFF;
                    11'h6AA : DATO <= 32'hFFFFFFFF;
                    11'h6AB : DATO <= 32'hFFFFFFFF;
                    11'h6AC : DATO <= 32'hFFFFFFFF;
                    11'h6AD : DATO <= 32'hFFFFFFFF;
                    11'h6AE : DATO <= 32'hFFFFFFFF;
                    11'h6AF : DATO <= 32'hFFFFFFFF;
                    11'h6B0 : DATO <= 32'hFFFFFFFF;
                    11'h6B1 : DATO <= 32'hFFFFFFFF;
                    11'h6B2 : DATO <= 32'hFFFFFFFF;
                    11'h6B3 : DATO <= 32'hFFFFFFFF;
                    11'h6B4 : DATO <= 32'hFFFFFFFF;
                    11'h6B5 : DATO <= 32'hFFFFFFFF;
                    11'h6B6 : DATO <= 32'hFFFFFFFF;
                    11'h6B7 : DATO <= 32'hFFFFFFFF;
                    11'h6B8 : DATO <= 32'hFFFFFFFF;
                    11'h6B9 : DATO <= 32'hFFFFFFFF;
                    11'h6BA : DATO <= 32'hFFFFFFFF;
                    11'h6BB : DATO <= 32'hFFFFFFFF;
                    11'h6BC : DATO <= 32'hFFFFFFFF;
                    11'h6BD : DATO <= 32'hFFFFFFFF;
                    11'h6BE : DATO <= 32'hFFFFFFFF;
                    11'h6BF : DATO <= 32'hFFFFFFFF;
                    11'h6C0 : DATO <= 32'hFFFFFFFF;
                    11'h6C1 : DATO <= 32'hFFFFFFFF;
                    11'h6C2 : DATO <= 32'hFFFFFFFF;
                    11'h6C3 : DATO <= 32'hFFFFFFFF;
                    11'h6C4 : DATO <= 32'hFFFFFFFF;
                    11'h6C5 : DATO <= 32'hFFFFFFFF;
                    11'h6C6 : DATO <= 32'hFFFFFFFF;
                    11'h6C7 : DATO <= 32'hFFFFFFFF;
                    11'h6C8 : DATO <= 32'hFFFFFFFF;
                    11'h6C9 : DATO <= 32'hFFFFFFFF;
                    11'h6CA : DATO <= 32'hFFFFFFFF;
                    11'h6CB : DATO <= 32'hFFFFFFFF;
                    11'h6CC : DATO <= 32'hFFFFFFFF;
                    11'h6CD : DATO <= 32'hFFFFFFFF;
                    11'h6CE : DATO <= 32'hFFFFFFFF;
                    11'h6CF : DATO <= 32'hFFFFFFFF;
                    11'h6D0 : DATO <= 32'hFFFFFFFF;
                    11'h6D1 : DATO <= 32'hFFFFFFFF;
                    11'h6D2 : DATO <= 32'hFFFFFFFF;
                    11'h6D3 : DATO <= 32'hFFFFFFFF;
                    11'h6D4 : DATO <= 32'hFFFFFFFF;
                    11'h6D5 : DATO <= 32'hFFFFFFFF;
                    11'h6D6 : DATO <= 32'hFFFFFFFF;
                    11'h6D7 : DATO <= 32'hFFFFFFFF;
                    11'h6D8 : DATO <= 32'hFFFFFFFF;
                    11'h6D9 : DATO <= 32'hFFFFFFFF;
                    11'h6DA : DATO <= 32'hFFFFFFFF;
                    11'h6DB : DATO <= 32'hFFFFFFFF;
                    11'h6DC : DATO <= 32'hFFFFFFFF;
                    11'h6DD : DATO <= 32'hFFFFFFFF;
                    11'h6DE : DATO <= 32'hFFFFFFFF;
                    11'h6DF : DATO <= 32'hFFFFFFFF;
                    11'h6E0 : DATO <= 32'hFFFFFFFF;
                    11'h6E1 : DATO <= 32'hFFFFFFFF;
                    11'h6E2 : DATO <= 32'hFFFFFFFF;
                    11'h6E3 : DATO <= 32'hFFFFFFFF;
                    11'h6E4 : DATO <= 32'hFFFFFFFF;
                    11'h6E5 : DATO <= 32'hFFFFFFFF;
                    11'h6E6 : DATO <= 32'hFFFFFFFF;
                    11'h6E7 : DATO <= 32'hFFFFFFFF;
                    11'h6E8 : DATO <= 32'hFFFFFFFF;
                    11'h6E9 : DATO <= 32'hFFFFFFFF;
                    11'h6EA : DATO <= 32'hFFFFFFFF;
                    11'h6EB : DATO <= 32'hFFFFFFFF;
                    11'h6EC : DATO <= 32'hFFFFFFFF;
                    11'h6ED : DATO <= 32'hFFFFFFFF;
                    11'h6EE : DATO <= 32'hFFFFFFFF;
                    11'h6EF : DATO <= 32'hFFFFFFFF;
                    11'h6F0 : DATO <= 32'hFFFFFFFF;
                    11'h6F1 : DATO <= 32'hFFFFFFFF;
                    11'h6F2 : DATO <= 32'hFFFFFFFF;
                    11'h6F3 : DATO <= 32'hFFFFFFFF;
                    11'h6F4 : DATO <= 32'hFFFFFFFF;
                    11'h6F5 : DATO <= 32'hFFFFFFFF;
                    11'h6F6 : DATO <= 32'hFFFFFFFF;
                    11'h6F7 : DATO <= 32'hFFFFFFFF;
                    11'h6F8 : DATO <= 32'hFFFFFFFF;
                    11'h6F9 : DATO <= 32'hFFFFFFFF;
                    11'h6FA : DATO <= 32'hFFFFFFFF;
                    11'h6FB : DATO <= 32'hFFFFFFFF;
                    11'h6FC : DATO <= 32'hFFFFFFFF;
                    11'h6FD : DATO <= 32'hFFFFFFFF;
                    11'h6FE : DATO <= 32'hFFFFFFFF;
                    11'h6FF : DATO <= 32'hFFFFFFFF;
                    11'h700 : DATO <= 32'hFFFFFFFF;
                    11'h701 : DATO <= 32'hFFFFFFFF;
                    11'h702 : DATO <= 32'hFFFFFFFF;
                    11'h703 : DATO <= 32'hFFFFFFFF;
                    11'h704 : DATO <= 32'hFFFFFFFF;
                    11'h705 : DATO <= 32'hFFFFFFFF;
                    11'h706 : DATO <= 32'hFFFFFFFF;
                    11'h707 : DATO <= 32'hFFFFFFFF;
                    11'h708 : DATO <= 32'hFFFFFFFF;
                    11'h709 : DATO <= 32'hFFFFFFFF;
                    11'h70A : DATO <= 32'hFFFFFFFF;
                    11'h70B : DATO <= 32'hFFFFFFFF;
                    11'h70C : DATO <= 32'hFFFFFFFF;
                    11'h70D : DATO <= 32'hFFFFFFFF;
                    11'h70E : DATO <= 32'hFFFFFFFF;
                    11'h70F : DATO <= 32'hFFFFFFFF;
                    11'h710 : DATO <= 32'hFFFFFFFF;
                    11'h711 : DATO <= 32'hFFFFFFFF;
                    11'h712 : DATO <= 32'hFFFFFFFF;
                    11'h713 : DATO <= 32'hFFFFFFFF;
                    11'h714 : DATO <= 32'hFFFFFFFF;
                    11'h715 : DATO <= 32'hFFFFFFFF;
                    11'h716 : DATO <= 32'hFFFFFFFF;
                    11'h717 : DATO <= 32'hFFFFFFFF;
                    11'h718 : DATO <= 32'hFFFFFFFF;
                    11'h719 : DATO <= 32'hFFFFFFFF;
                    11'h71A : DATO <= 32'hFFFFFFFF;
                    11'h71B : DATO <= 32'hFFFFFFFF;
                    11'h71C : DATO <= 32'hFFFFFFFF;
                    11'h71D : DATO <= 32'hFFFFFFFF;
                    11'h71E : DATO <= 32'hFFFFFFFF;
                    11'h71F : DATO <= 32'hFFFFFFFF;
                    11'h720 : DATO <= 32'hFFFFFFFF;
                    11'h721 : DATO <= 32'hFFFFFFFF;
                    11'h722 : DATO <= 32'hFFFFFFFF;
                    11'h723 : DATO <= 32'hFFFFFFFF;
                    11'h724 : DATO <= 32'hFFFFFFFF;
                    11'h725 : DATO <= 32'hFFFFFFFF;
                    11'h726 : DATO <= 32'hFFFFFFFF;
                    11'h727 : DATO <= 32'hFFFFFFFF;
                    11'h728 : DATO <= 32'hFFFFFFFF;
                    11'h729 : DATO <= 32'hFFFFFFFF;
                    11'h72A : DATO <= 32'hFFFFFFFF;
                    11'h72B : DATO <= 32'hFFFFFFFF;
                    11'h72C : DATO <= 32'hFFFFFFFF;
                    11'h72D : DATO <= 32'hFFFFFFFF;
                    11'h72E : DATO <= 32'hFFFFFFFF;
                    11'h72F : DATO <= 32'hFFFFFFFF;
                    11'h730 : DATO <= 32'hFFFFFFFF;
                    11'h731 : DATO <= 32'hFFFFFFFF;
                    11'h732 : DATO <= 32'hFFFFFFFF;
                    11'h733 : DATO <= 32'hFFFFFFFF;
                    11'h734 : DATO <= 32'hFFFFFFFF;
                    11'h735 : DATO <= 32'hFFFFFFFF;
                    11'h736 : DATO <= 32'hFFFFFFFF;
                    11'h737 : DATO <= 32'hFFFFFFFF;
                    11'h738 : DATO <= 32'hFFFFFFFF;
                    11'h739 : DATO <= 32'hFFFFFFFF;
                    11'h73A : DATO <= 32'hFFFFFFFF;
                    11'h73B : DATO <= 32'hFFFFFFFF;
                    11'h73C : DATO <= 32'hFFFFFFFF;
                    11'h73D : DATO <= 32'hFFFFFFFF;
                    11'h73E : DATO <= 32'hFFFFFFFF;
                    11'h73F : DATO <= 32'hFFFFFFFF;
                    11'h740 : DATO <= 32'hFFFFFFFF;
                    11'h741 : DATO <= 32'hFFFFFFFF;
                    11'h742 : DATO <= 32'hFFFFFFFF;
                    11'h743 : DATO <= 32'hFFFFFFFF;
                    11'h744 : DATO <= 32'hFFFFFFFF;
                    11'h745 : DATO <= 32'hFFFFFFFF;
                    11'h746 : DATO <= 32'hFFFFFFFF;
                    11'h747 : DATO <= 32'hFFFFFFFF;
                    11'h748 : DATO <= 32'hFFFFFFFF;
                    11'h749 : DATO <= 32'hFFFFFFFF;
                    11'h74A : DATO <= 32'hFFFFFFFF;
                    11'h74B : DATO <= 32'hFFFFFFFF;
                    11'h74C : DATO <= 32'hFFFFFFFF;
                    11'h74D : DATO <= 32'hFFFFFFFF;
                    11'h74E : DATO <= 32'hFFFFFFFF;
                    11'h74F : DATO <= 32'hFFFFFFFF;
                    11'h750 : DATO <= 32'hFFFFFFFF;
                    11'h751 : DATO <= 32'hFFFFFFFF;
                    11'h752 : DATO <= 32'hFFFFFFFF;
                    11'h753 : DATO <= 32'hFFFFFFFF;
                    11'h754 : DATO <= 32'hFFFFFFFF;
                    11'h755 : DATO <= 32'hFFFFFFFF;
                    11'h756 : DATO <= 32'hFFFFFFFF;
                    11'h757 : DATO <= 32'hFFFFFFFF;
                    11'h758 : DATO <= 32'hFFFFFFFF;
                    11'h759 : DATO <= 32'hFFFFFFFF;
                    11'h75A : DATO <= 32'hFFFFFFFF;
                    11'h75B : DATO <= 32'hFFFFFFFF;
                    11'h75C : DATO <= 32'hFFFFFFFF;
                    11'h75D : DATO <= 32'hFFFFFFFF;
                    11'h75E : DATO <= 32'hFFFFFFFF;
                    11'h75F : DATO <= 32'hFFFFFFFF;
                    11'h760 : DATO <= 32'hFFFFFFFF;
                    11'h761 : DATO <= 32'hFFFFFFFF;
                    11'h762 : DATO <= 32'hFFFFFFFF;
                    11'h763 : DATO <= 32'hFFFFFFFF;
                    11'h764 : DATO <= 32'hFFFFFFFF;
                    11'h765 : DATO <= 32'hFFFFFFFF;
                    11'h766 : DATO <= 32'hFFFFFFFF;
                    11'h767 : DATO <= 32'hFFFFFFFF;
                    11'h768 : DATO <= 32'hFFFFFFFF;
                    11'h769 : DATO <= 32'hFFFFFFFF;
                    11'h76A : DATO <= 32'hFFFFFFFF;
                    11'h76B : DATO <= 32'hFFFFFFFF;
                    11'h76C : DATO <= 32'hFFFFFFFF;
                    11'h76D : DATO <= 32'hFFFFFFFF;
                    11'h76E : DATO <= 32'hFFFFFFFF;
                    11'h76F : DATO <= 32'hFFFFFFFF;
                    11'h770 : DATO <= 32'hFFFFFFFF;
                    11'h771 : DATO <= 32'hFFFFFFFF;
                    11'h772 : DATO <= 32'hFFFFFFFF;
                    11'h773 : DATO <= 32'hFFFFFFFF;
                    11'h774 : DATO <= 32'hFFFFFFFF;
                    11'h775 : DATO <= 32'hFFFFFFFF;
                    11'h776 : DATO <= 32'hFFFFFFFF;
                    11'h777 : DATO <= 32'hFFFFFFFF;
                    11'h778 : DATO <= 32'hFFFFFFFF;
                    11'h779 : DATO <= 32'hFFFFFFFF;
                    11'h77A : DATO <= 32'hFFFFFFFF;
                    11'h77B : DATO <= 32'hFFFFFFFF;
                    11'h77C : DATO <= 32'hFFFFFFFF;
                    11'h77D : DATO <= 32'hFFFFFFFF;
                    11'h77E : DATO <= 32'hFFFFFFFF;
                    11'h77F : DATO <= 32'hFFFFFFFF;
                    11'h780 : DATO <= 32'hFFFFFFFF;
                    11'h781 : DATO <= 32'hFFFFFFFF;
                    11'h782 : DATO <= 32'hFFFFFFFF;
                    11'h783 : DATO <= 32'hFFFFFFFF;
                    11'h784 : DATO <= 32'hFFFFFFFF;
                    11'h785 : DATO <= 32'hFFFFFFFF;
                    11'h786 : DATO <= 32'hFFFFFFFF;
                    11'h787 : DATO <= 32'hFFFFFFFF;
                    11'h788 : DATO <= 32'hFFFFFFFF;
                    11'h789 : DATO <= 32'hFFFFFFFF;
                    11'h78A : DATO <= 32'hFFFFFFFF;
                    11'h78B : DATO <= 32'hFFFFFFFF;
                    11'h78C : DATO <= 32'hFFFFFFFF;
                    11'h78D : DATO <= 32'hFFFFFFFF;
                    11'h78E : DATO <= 32'hFFFFFFFF;
                    11'h78F : DATO <= 32'hFFFFFFFF;
                    11'h790 : DATO <= 32'hFFFFFFFF;
                    11'h791 : DATO <= 32'hFFFFFFFF;
                    11'h792 : DATO <= 32'hFFFFFFFF;
                    11'h793 : DATO <= 32'hFFFFFFFF;
                    11'h794 : DATO <= 32'hFFFFFFFF;
                    11'h795 : DATO <= 32'hFFFFFFFF;
                    11'h796 : DATO <= 32'hFFFFFFFF;
                    11'h797 : DATO <= 32'hFFFFFFFF;
                    11'h798 : DATO <= 32'hFFFFFFFF;
                    11'h799 : DATO <= 32'hFFFFFFFF;
                    11'h79A : DATO <= 32'hFFFFFFFF;
                    11'h79B : DATO <= 32'hFFFFFFFF;
                    11'h79C : DATO <= 32'hFFFFFFFF;
                    11'h79D : DATO <= 32'hFFFFFFFF;
                    11'h79E : DATO <= 32'hFFFFFFFF;
                    11'h79F : DATO <= 32'hFFFFFFFF;
                    11'h7A0 : DATO <= 32'hFFFFFFFF;
                    11'h7A1 : DATO <= 32'hFFFFFFFF;
                    11'h7A2 : DATO <= 32'hFFFFFFFF;
                    11'h7A3 : DATO <= 32'hFFFFFFFF;
                    11'h7A4 : DATO <= 32'hFFFFFFFF;
                    11'h7A5 : DATO <= 32'hFFFFFFFF;
                    11'h7A6 : DATO <= 32'hFFFFFFFF;
                    11'h7A7 : DATO <= 32'hFFFFFFFF;
                    11'h7A8 : DATO <= 32'hFFFFFFFF;
                    11'h7A9 : DATO <= 32'hFFFFFFFF;
                    11'h7AA : DATO <= 32'hFFFFFFFF;
                    11'h7AB : DATO <= 32'hFFFFFFFF;
                    11'h7AC : DATO <= 32'hFFFFFFFF;
                    11'h7AD : DATO <= 32'hFFFFFFFF;
                    11'h7AE : DATO <= 32'hFFFFFFFF;
                    11'h7AF : DATO <= 32'hFFFFFFFF;
                    11'h7B0 : DATO <= 32'hFFFFFFFF;
                    11'h7B1 : DATO <= 32'hFFFFFFFF;
                    11'h7B2 : DATO <= 32'hFFFFFFFF;
                    11'h7B3 : DATO <= 32'hFFFFFFFF;
                    11'h7B4 : DATO <= 32'hFFFFFFFF;
                    11'h7B5 : DATO <= 32'hFFFFFFFF;
                    11'h7B6 : DATO <= 32'hFFFFFFFF;
                    11'h7B7 : DATO <= 32'hFFFFFFFF;
                    11'h7B8 : DATO <= 32'hFFFFFFFF;
                    11'h7B9 : DATO <= 32'hFFFFFFFF;
                    11'h7BA : DATO <= 32'hFFFFFFFF;
                    11'h7BB : DATO <= 32'hFFFFFFFF;
                    11'h7BC : DATO <= 32'hFFFFFFFF;
                    11'h7BD : DATO <= 32'hFFFFFFFF;
                    11'h7BE : DATO <= 32'hFFFFFFFF;
                    11'h7BF : DATO <= 32'hFFFFFFFF;
                    11'h7C0 : DATO <= 32'hFFFFFFFF;
                    11'h7C1 : DATO <= 32'hFFFFFFFF;
                    11'h7C2 : DATO <= 32'hFFFFFFFF;
                    11'h7C3 : DATO <= 32'hFFFFFFFF;
                    11'h7C4 : DATO <= 32'hFFFFFFFF;
                    11'h7C5 : DATO <= 32'hFFFFFFFF;
                    11'h7C6 : DATO <= 32'hFFFFFFFF;
                    11'h7C7 : DATO <= 32'hFFFFFFFF;
                    11'h7C8 : DATO <= 32'hFFFFFFFF;
                    11'h7C9 : DATO <= 32'hFFFFFFFF;
                    11'h7CA : DATO <= 32'hFFFFFFFF;
                    11'h7CB : DATO <= 32'hFFFFFFFF;
                    11'h7CC : DATO <= 32'hFFFFFFFF;
                    11'h7CD : DATO <= 32'hFFFFFFFF;
                    11'h7CE : DATO <= 32'hFFFFFFFF;
                    11'h7CF : DATO <= 32'hFFFFFFFF;
                    11'h7D0 : DATO <= 32'hFFFFFFFF;
                    11'h7D1 : DATO <= 32'hFFFFFFFF;
                    11'h7D2 : DATO <= 32'hFFFFFFFF;
                    11'h7D3 : DATO <= 32'hFFFFFFFF;
                    11'h7D4 : DATO <= 32'hFFFFFFFF;
                    11'h7D5 : DATO <= 32'hFFFFFFFF;
                    11'h7D6 : DATO <= 32'hFFFFFFFF;
                    11'h7D7 : DATO <= 32'hFFFFFFFF;
                    11'h7D8 : DATO <= 32'hFFFFFFFF;
                    11'h7D9 : DATO <= 32'hFFFFFFFF;
                    11'h7DA : DATO <= 32'hFFFFFFFF;
                    11'h7DB : DATO <= 32'hFFFFFFFF;
                    11'h7DC : DATO <= 32'hFFFFFFFF;
                    11'h7DD : DATO <= 32'hFFFFFFFF;
                    11'h7DE : DATO <= 32'hFFFFFFFF;
                    11'h7DF : DATO <= 32'hFFFFFFFF;
                    11'h7E0 : DATO <= 32'hFFFFFFFF;
                    11'h7E1 : DATO <= 32'hFFFFFFFF;
                    11'h7E2 : DATO <= 32'hFFFFFFFF;
                    11'h7E3 : DATO <= 32'hFFFFFFFF;
                    11'h7E4 : DATO <= 32'hFFFFFFFF;
                    11'h7E5 : DATO <= 32'hFFFFFFFF;
                    11'h7E6 : DATO <= 32'hFFFFFFFF;
                    11'h7E7 : DATO <= 32'hFFFFFFFF;
                    11'h7E8 : DATO <= 32'hFFFFFFFF;
                    11'h7E9 : DATO <= 32'hFFFFFFFF;
                    11'h7EA : DATO <= 32'hFFFFFFFF;
                    11'h7EB : DATO <= 32'hFFFFFFFF;
                    11'h7EC : DATO <= 32'hFFFFFFFF;
                    11'h7ED : DATO <= 32'hFFFFFFFF;
                    11'h7EE : DATO <= 32'hFFFFFFFF;
                    11'h7EF : DATO <= 32'hFFFFFFFF;
                    11'h7F0 : DATO <= 32'hFFFFFFFF;
                    11'h7F1 : DATO <= 32'hFFFFFFFF;
                    11'h7F2 : DATO <= 32'hFFFFFFFF;
                    11'h7F3 : DATO <= 32'hFFFFFFFF;
                    11'h7F4 : DATO <= 32'hFFFFFFFF;
                    11'h7F5 : DATO <= 32'hFFFFFFFF;
                    11'h7F6 : DATO <= 32'hFFFFFFFF;
                    11'h7F7 : DATO <= 32'hFFFFFFFF;
                    11'h7F8 : DATO <= 32'hFFFFFFFF;
                    11'h7F9 : DATO <= 32'hFFFFFFFF;
                    11'h7FA : DATO <= 32'hFFFFFFFF;
                    11'h7FB : DATO <= 32'hFFFFFFFF;
                    11'h7FC : DATO <= 32'hFFFFFFFF;
                    11'h7FD : DATO <= 32'hFFFFFFFF;
                    11'h7FE : DATO <= 32'hFFFFFFFF;
                    11'h7FF : DATO <= 32'hFFFFFFFF;
                    default : DATO <= 32'hxxxxxxxx;
                endcase
            end
    end
endmodule
