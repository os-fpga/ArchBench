//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for physical tile: io_right_top]
//	Author: Xifan TANG
//	Organization: University of Utah
//-------------------------------------------
//----- Time scale -----
`timescale 1ns / 1ps

// ----- BEGIN Grid Verilog module: grid_io_right_top -----
//----- Default net type -----
`default_nettype wire

// ----- Verilog module for grid_io_right_top -----
module grid_io_right_top(global_reset,
                         scan_mode,
                         scan_enable,
                         config_enable,
                         prog_clock,
                         gfpga_pad_RS_PREIO_A2F,
                         gfpga_pad_RS_PREIO_F2A,
                         gfpga_pad_RS_PREIO_SOC_CLK,
                         top_width_0_height_0_subtile_14__pin_f2a_i_0_,
                         top_width_0_height_0_subtile_15__pin_f2a_i_0_,
                         top_width_0_height_0_subtile_16__pin_f2a_i_0_,
                         top_width_0_height_0_subtile_17__pin_f2a_i_0_,
                         top_width_0_height_0_subtile_18__pin_f2a_i_0_,
                         top_width_0_height_0_subtile_19__pin_f2a_i_0_,
                         top_width_0_height_0_subtile_20__pin_f2a_i_0_,
                         top_width_0_height_0_subtile_21__pin_f2a_i_0_,
                         top_width_0_height_0_subtile_22__pin_f2a_i_0_,
                         top_width_0_height_0_subtile_23__pin_f2a_i_0_,
                         top_width_0_height_0_subtile_24__pin_f2a_i_0_,
                         top_width_0_height_0_subtile_25__pin_f2a_i_0_,
                         top_width_0_height_0_subtile_26__pin_f2a_i_0_,
                         top_width_0_height_0_subtile_27__pin_f2a_i_0_,
                         top_width_0_height_0_subtile_28__pin_f2a_i_0_,
                         top_width_0_height_0_subtile_29__pin_f2a_i_0_,
                         top_width_0_height_0_subtile_30__pin_f2a_i_0_,
                         top_width_0_height_0_subtile_31__pin_f2a_i_0_,
                         top_width_0_height_0_subtile_32__pin_f2a_i_0_,
                         top_width_0_height_0_subtile_33__pin_f2a_i_0_,
                         top_width_0_height_0_subtile_34__pin_f2a_i_0_,
                         top_width_0_height_0_subtile_35__pin_f2a_i_0_,
                         top_width_0_height_0_subtile_36__pin_f2a_i_0_,
                         top_width_0_height_0_subtile_37__pin_f2a_i_0_,
                         top_width_0_height_0_subtile_38__pin_f2a_i_0_,
                         top_width_0_height_0_subtile_39__pin_f2a_i_0_,
                         top_width_0_height_0_subtile_40__pin_f2a_i_0_,
                         top_width_0_height_0_subtile_41__pin_f2a_i_0_,
                         top_width_0_height_0_subtile_42__pin_f2a_i_0_,
                         top_width_0_height_0_subtile_43__pin_f2a_i_0_,
                         top_width_0_height_0_subtile_44__pin_f2a_i_0_,
                         top_width_0_height_0_subtile_45__pin_f2a_i_0_,
                         top_width_0_height_0_subtile_46__pin_f2a_i_0_,
                         top_width_0_height_0_subtile_47__pin_f2a_i_0_,
                         top_width_0_height_0_subtile_48__pin_f2a_i_0_,
                         top_width_0_height_0_subtile_49__pin_f2a_i_0_,
                         top_width_0_height_0_subtile_50__pin_f2a_i_0_,
                         top_width_0_height_0_subtile_51__pin_f2a_i_0_,
                         top_width_0_height_0_subtile_52__pin_f2a_i_0_,
                         top_width_0_height_0_subtile_53__pin_f2a_i_0_,
                         top_width_0_height_0_subtile_54__pin_f2a_i_0_,
                         top_width_0_height_0_subtile_55__pin_f2a_i_0_,
                         top_width_0_height_0_subtile_56__pin_f2a_i_0_,
                         top_width_0_height_0_subtile_57__pin_f2a_i_0_,
                         top_width_0_height_0_subtile_58__pin_f2a_i_0_,
                         top_width_0_height_0_subtile_59__pin_f2a_i_0_,
                         right_width_0_height_0_subtile_0__pin_f2a_i_0_,
                         right_width_0_height_0_subtile_1__pin_f2a_i_0_,
                         right_width_0_height_0_subtile_2__pin_f2a_i_0_,
                         right_width_0_height_0_subtile_3__pin_f2a_i_0_,
                         right_width_0_height_0_subtile_4__pin_f2a_i_0_,
                         right_width_0_height_0_subtile_5__pin_f2a_i_0_,
                         right_width_0_height_0_subtile_6__pin_f2a_i_0_,
                         right_width_0_height_0_subtile_7__pin_f2a_i_0_,
                         right_width_0_height_0_subtile_8__pin_f2a_i_0_,
                         right_width_0_height_0_subtile_9__pin_f2a_i_0_,
                         right_width_0_height_0_subtile_10__pin_f2a_i_0_,
                         right_width_0_height_0_subtile_11__pin_f2a_i_0_,
                         right_width_0_height_0_subtile_12__pin_f2a_i_0_,
                         right_width_0_height_0_subtile_13__pin_f2a_i_0_,
                         bottom_width_0_height_0_subtile_0__pin_clk_0_,
                         bottom_width_0_height_0_subtile_0__pin_clk_1_,
                         bottom_width_0_height_0_subtile_0__pin_clk_2_,
                         bottom_width_0_height_0_subtile_0__pin_clk_3_,
                         bottom_width_0_height_0_subtile_0__pin_clk_4_,
                         bottom_width_0_height_0_subtile_0__pin_clk_5_,
                         bottom_width_0_height_0_subtile_0__pin_clk_6_,
                         bottom_width_0_height_0_subtile_0__pin_clk_7_,
                         bottom_width_0_height_0_subtile_0__pin_clk_8_,
                         bottom_width_0_height_0_subtile_0__pin_clk_9_,
                         bottom_width_0_height_0_subtile_0__pin_clk_10_,
                         bottom_width_0_height_0_subtile_0__pin_clk_11_,
                         bottom_width_0_height_0_subtile_0__pin_clk_12_,
                         bottom_width_0_height_0_subtile_0__pin_clk_13_,
                         bottom_width_0_height_0_subtile_0__pin_clk_14_,
                         bottom_width_0_height_0_subtile_0__pin_clk_15_,
                         bottom_width_0_height_0_subtile_1__pin_clk_0_,
                         bottom_width_0_height_0_subtile_1__pin_clk_1_,
                         bottom_width_0_height_0_subtile_1__pin_clk_2_,
                         bottom_width_0_height_0_subtile_1__pin_clk_3_,
                         bottom_width_0_height_0_subtile_1__pin_clk_4_,
                         bottom_width_0_height_0_subtile_1__pin_clk_5_,
                         bottom_width_0_height_0_subtile_1__pin_clk_6_,
                         bottom_width_0_height_0_subtile_1__pin_clk_7_,
                         bottom_width_0_height_0_subtile_1__pin_clk_8_,
                         bottom_width_0_height_0_subtile_1__pin_clk_9_,
                         bottom_width_0_height_0_subtile_1__pin_clk_10_,
                         bottom_width_0_height_0_subtile_1__pin_clk_11_,
                         bottom_width_0_height_0_subtile_1__pin_clk_12_,
                         bottom_width_0_height_0_subtile_1__pin_clk_13_,
                         bottom_width_0_height_0_subtile_1__pin_clk_14_,
                         bottom_width_0_height_0_subtile_1__pin_clk_15_,
                         bottom_width_0_height_0_subtile_2__pin_clk_0_,
                         bottom_width_0_height_0_subtile_2__pin_clk_1_,
                         bottom_width_0_height_0_subtile_2__pin_clk_2_,
                         bottom_width_0_height_0_subtile_2__pin_clk_3_,
                         bottom_width_0_height_0_subtile_2__pin_clk_4_,
                         bottom_width_0_height_0_subtile_2__pin_clk_5_,
                         bottom_width_0_height_0_subtile_2__pin_clk_6_,
                         bottom_width_0_height_0_subtile_2__pin_clk_7_,
                         bottom_width_0_height_0_subtile_2__pin_clk_8_,
                         bottom_width_0_height_0_subtile_2__pin_clk_9_,
                         bottom_width_0_height_0_subtile_2__pin_clk_10_,
                         bottom_width_0_height_0_subtile_2__pin_clk_11_,
                         bottom_width_0_height_0_subtile_2__pin_clk_12_,
                         bottom_width_0_height_0_subtile_2__pin_clk_13_,
                         bottom_width_0_height_0_subtile_2__pin_clk_14_,
                         bottom_width_0_height_0_subtile_2__pin_clk_15_,
                         bottom_width_0_height_0_subtile_3__pin_clk_0_,
                         bottom_width_0_height_0_subtile_3__pin_clk_1_,
                         bottom_width_0_height_0_subtile_3__pin_clk_2_,
                         bottom_width_0_height_0_subtile_3__pin_clk_3_,
                         bottom_width_0_height_0_subtile_3__pin_clk_4_,
                         bottom_width_0_height_0_subtile_3__pin_clk_5_,
                         bottom_width_0_height_0_subtile_3__pin_clk_6_,
                         bottom_width_0_height_0_subtile_3__pin_clk_7_,
                         bottom_width_0_height_0_subtile_3__pin_clk_8_,
                         bottom_width_0_height_0_subtile_3__pin_clk_9_,
                         bottom_width_0_height_0_subtile_3__pin_clk_10_,
                         bottom_width_0_height_0_subtile_3__pin_clk_11_,
                         bottom_width_0_height_0_subtile_3__pin_clk_12_,
                         bottom_width_0_height_0_subtile_3__pin_clk_13_,
                         bottom_width_0_height_0_subtile_3__pin_clk_14_,
                         bottom_width_0_height_0_subtile_3__pin_clk_15_,
                         bottom_width_0_height_0_subtile_4__pin_clk_0_,
                         bottom_width_0_height_0_subtile_4__pin_clk_1_,
                         bottom_width_0_height_0_subtile_4__pin_clk_2_,
                         bottom_width_0_height_0_subtile_4__pin_clk_3_,
                         bottom_width_0_height_0_subtile_4__pin_clk_4_,
                         bottom_width_0_height_0_subtile_4__pin_clk_5_,
                         bottom_width_0_height_0_subtile_4__pin_clk_6_,
                         bottom_width_0_height_0_subtile_4__pin_clk_7_,
                         bottom_width_0_height_0_subtile_4__pin_clk_8_,
                         bottom_width_0_height_0_subtile_4__pin_clk_9_,
                         bottom_width_0_height_0_subtile_4__pin_clk_10_,
                         bottom_width_0_height_0_subtile_4__pin_clk_11_,
                         bottom_width_0_height_0_subtile_4__pin_clk_12_,
                         bottom_width_0_height_0_subtile_4__pin_clk_13_,
                         bottom_width_0_height_0_subtile_4__pin_clk_14_,
                         bottom_width_0_height_0_subtile_4__pin_clk_15_,
                         bottom_width_0_height_0_subtile_5__pin_clk_0_,
                         bottom_width_0_height_0_subtile_5__pin_clk_1_,
                         bottom_width_0_height_0_subtile_5__pin_clk_2_,
                         bottom_width_0_height_0_subtile_5__pin_clk_3_,
                         bottom_width_0_height_0_subtile_5__pin_clk_4_,
                         bottom_width_0_height_0_subtile_5__pin_clk_5_,
                         bottom_width_0_height_0_subtile_5__pin_clk_6_,
                         bottom_width_0_height_0_subtile_5__pin_clk_7_,
                         bottom_width_0_height_0_subtile_5__pin_clk_8_,
                         bottom_width_0_height_0_subtile_5__pin_clk_9_,
                         bottom_width_0_height_0_subtile_5__pin_clk_10_,
                         bottom_width_0_height_0_subtile_5__pin_clk_11_,
                         bottom_width_0_height_0_subtile_5__pin_clk_12_,
                         bottom_width_0_height_0_subtile_5__pin_clk_13_,
                         bottom_width_0_height_0_subtile_5__pin_clk_14_,
                         bottom_width_0_height_0_subtile_5__pin_clk_15_,
                         bottom_width_0_height_0_subtile_6__pin_clk_0_,
                         bottom_width_0_height_0_subtile_6__pin_clk_1_,
                         bottom_width_0_height_0_subtile_6__pin_clk_2_,
                         bottom_width_0_height_0_subtile_6__pin_clk_3_,
                         bottom_width_0_height_0_subtile_6__pin_clk_4_,
                         bottom_width_0_height_0_subtile_6__pin_clk_5_,
                         bottom_width_0_height_0_subtile_6__pin_clk_6_,
                         bottom_width_0_height_0_subtile_6__pin_clk_7_,
                         bottom_width_0_height_0_subtile_6__pin_clk_8_,
                         bottom_width_0_height_0_subtile_6__pin_clk_9_,
                         bottom_width_0_height_0_subtile_6__pin_clk_10_,
                         bottom_width_0_height_0_subtile_6__pin_clk_11_,
                         bottom_width_0_height_0_subtile_6__pin_clk_12_,
                         bottom_width_0_height_0_subtile_6__pin_clk_13_,
                         bottom_width_0_height_0_subtile_6__pin_clk_14_,
                         bottom_width_0_height_0_subtile_6__pin_clk_15_,
                         bottom_width_0_height_0_subtile_7__pin_clk_0_,
                         bottom_width_0_height_0_subtile_7__pin_clk_1_,
                         bottom_width_0_height_0_subtile_7__pin_clk_2_,
                         bottom_width_0_height_0_subtile_7__pin_clk_3_,
                         bottom_width_0_height_0_subtile_7__pin_clk_4_,
                         bottom_width_0_height_0_subtile_7__pin_clk_5_,
                         bottom_width_0_height_0_subtile_7__pin_clk_6_,
                         bottom_width_0_height_0_subtile_7__pin_clk_7_,
                         bottom_width_0_height_0_subtile_7__pin_clk_8_,
                         bottom_width_0_height_0_subtile_7__pin_clk_9_,
                         bottom_width_0_height_0_subtile_7__pin_clk_10_,
                         bottom_width_0_height_0_subtile_7__pin_clk_11_,
                         bottom_width_0_height_0_subtile_7__pin_clk_12_,
                         bottom_width_0_height_0_subtile_7__pin_clk_13_,
                         bottom_width_0_height_0_subtile_7__pin_clk_14_,
                         bottom_width_0_height_0_subtile_7__pin_clk_15_,
                         bottom_width_0_height_0_subtile_8__pin_clk_0_,
                         bottom_width_0_height_0_subtile_8__pin_clk_1_,
                         bottom_width_0_height_0_subtile_8__pin_clk_2_,
                         bottom_width_0_height_0_subtile_8__pin_clk_3_,
                         bottom_width_0_height_0_subtile_8__pin_clk_4_,
                         bottom_width_0_height_0_subtile_8__pin_clk_5_,
                         bottom_width_0_height_0_subtile_8__pin_clk_6_,
                         bottom_width_0_height_0_subtile_8__pin_clk_7_,
                         bottom_width_0_height_0_subtile_8__pin_clk_8_,
                         bottom_width_0_height_0_subtile_8__pin_clk_9_,
                         bottom_width_0_height_0_subtile_8__pin_clk_10_,
                         bottom_width_0_height_0_subtile_8__pin_clk_11_,
                         bottom_width_0_height_0_subtile_8__pin_clk_12_,
                         bottom_width_0_height_0_subtile_8__pin_clk_13_,
                         bottom_width_0_height_0_subtile_8__pin_clk_14_,
                         bottom_width_0_height_0_subtile_8__pin_clk_15_,
                         bottom_width_0_height_0_subtile_9__pin_clk_0_,
                         bottom_width_0_height_0_subtile_9__pin_clk_1_,
                         bottom_width_0_height_0_subtile_9__pin_clk_2_,
                         bottom_width_0_height_0_subtile_9__pin_clk_3_,
                         bottom_width_0_height_0_subtile_9__pin_clk_4_,
                         bottom_width_0_height_0_subtile_9__pin_clk_5_,
                         bottom_width_0_height_0_subtile_9__pin_clk_6_,
                         bottom_width_0_height_0_subtile_9__pin_clk_7_,
                         bottom_width_0_height_0_subtile_9__pin_clk_8_,
                         bottom_width_0_height_0_subtile_9__pin_clk_9_,
                         bottom_width_0_height_0_subtile_9__pin_clk_10_,
                         bottom_width_0_height_0_subtile_9__pin_clk_11_,
                         bottom_width_0_height_0_subtile_9__pin_clk_12_,
                         bottom_width_0_height_0_subtile_9__pin_clk_13_,
                         bottom_width_0_height_0_subtile_9__pin_clk_14_,
                         bottom_width_0_height_0_subtile_9__pin_clk_15_,
                         bottom_width_0_height_0_subtile_10__pin_clk_0_,
                         bottom_width_0_height_0_subtile_10__pin_clk_1_,
                         bottom_width_0_height_0_subtile_10__pin_clk_2_,
                         bottom_width_0_height_0_subtile_10__pin_clk_3_,
                         bottom_width_0_height_0_subtile_10__pin_clk_4_,
                         bottom_width_0_height_0_subtile_10__pin_clk_5_,
                         bottom_width_0_height_0_subtile_10__pin_clk_6_,
                         bottom_width_0_height_0_subtile_10__pin_clk_7_,
                         bottom_width_0_height_0_subtile_10__pin_clk_8_,
                         bottom_width_0_height_0_subtile_10__pin_clk_9_,
                         bottom_width_0_height_0_subtile_10__pin_clk_10_,
                         bottom_width_0_height_0_subtile_10__pin_clk_11_,
                         bottom_width_0_height_0_subtile_10__pin_clk_12_,
                         bottom_width_0_height_0_subtile_10__pin_clk_13_,
                         bottom_width_0_height_0_subtile_10__pin_clk_14_,
                         bottom_width_0_height_0_subtile_10__pin_clk_15_,
                         bottom_width_0_height_0_subtile_11__pin_clk_0_,
                         bottom_width_0_height_0_subtile_11__pin_clk_1_,
                         bottom_width_0_height_0_subtile_11__pin_clk_2_,
                         bottom_width_0_height_0_subtile_11__pin_clk_3_,
                         bottom_width_0_height_0_subtile_11__pin_clk_4_,
                         bottom_width_0_height_0_subtile_11__pin_clk_5_,
                         bottom_width_0_height_0_subtile_11__pin_clk_6_,
                         bottom_width_0_height_0_subtile_11__pin_clk_7_,
                         bottom_width_0_height_0_subtile_11__pin_clk_8_,
                         bottom_width_0_height_0_subtile_11__pin_clk_9_,
                         bottom_width_0_height_0_subtile_11__pin_clk_10_,
                         bottom_width_0_height_0_subtile_11__pin_clk_11_,
                         bottom_width_0_height_0_subtile_11__pin_clk_12_,
                         bottom_width_0_height_0_subtile_11__pin_clk_13_,
                         bottom_width_0_height_0_subtile_11__pin_clk_14_,
                         bottom_width_0_height_0_subtile_11__pin_clk_15_,
                         bottom_width_0_height_0_subtile_12__pin_clk_0_,
                         bottom_width_0_height_0_subtile_12__pin_clk_1_,
                         bottom_width_0_height_0_subtile_12__pin_clk_2_,
                         bottom_width_0_height_0_subtile_12__pin_clk_3_,
                         bottom_width_0_height_0_subtile_12__pin_clk_4_,
                         bottom_width_0_height_0_subtile_12__pin_clk_5_,
                         bottom_width_0_height_0_subtile_12__pin_clk_6_,
                         bottom_width_0_height_0_subtile_12__pin_clk_7_,
                         bottom_width_0_height_0_subtile_12__pin_clk_8_,
                         bottom_width_0_height_0_subtile_12__pin_clk_9_,
                         bottom_width_0_height_0_subtile_12__pin_clk_10_,
                         bottom_width_0_height_0_subtile_12__pin_clk_11_,
                         bottom_width_0_height_0_subtile_12__pin_clk_12_,
                         bottom_width_0_height_0_subtile_12__pin_clk_13_,
                         bottom_width_0_height_0_subtile_12__pin_clk_14_,
                         bottom_width_0_height_0_subtile_12__pin_clk_15_,
                         bottom_width_0_height_0_subtile_13__pin_clk_0_,
                         bottom_width_0_height_0_subtile_13__pin_clk_1_,
                         bottom_width_0_height_0_subtile_13__pin_clk_2_,
                         bottom_width_0_height_0_subtile_13__pin_clk_3_,
                         bottom_width_0_height_0_subtile_13__pin_clk_4_,
                         bottom_width_0_height_0_subtile_13__pin_clk_5_,
                         bottom_width_0_height_0_subtile_13__pin_clk_6_,
                         bottom_width_0_height_0_subtile_13__pin_clk_7_,
                         bottom_width_0_height_0_subtile_13__pin_clk_8_,
                         bottom_width_0_height_0_subtile_13__pin_clk_9_,
                         bottom_width_0_height_0_subtile_13__pin_clk_10_,
                         bottom_width_0_height_0_subtile_13__pin_clk_11_,
                         bottom_width_0_height_0_subtile_13__pin_clk_12_,
                         bottom_width_0_height_0_subtile_13__pin_clk_13_,
                         bottom_width_0_height_0_subtile_13__pin_clk_14_,
                         bottom_width_0_height_0_subtile_13__pin_clk_15_,
                         bottom_width_0_height_0_subtile_14__pin_clk_0_,
                         bottom_width_0_height_0_subtile_14__pin_clk_1_,
                         bottom_width_0_height_0_subtile_14__pin_clk_2_,
                         bottom_width_0_height_0_subtile_14__pin_clk_3_,
                         bottom_width_0_height_0_subtile_14__pin_clk_4_,
                         bottom_width_0_height_0_subtile_14__pin_clk_5_,
                         bottom_width_0_height_0_subtile_14__pin_clk_6_,
                         bottom_width_0_height_0_subtile_14__pin_clk_7_,
                         bottom_width_0_height_0_subtile_14__pin_clk_8_,
                         bottom_width_0_height_0_subtile_14__pin_clk_9_,
                         bottom_width_0_height_0_subtile_14__pin_clk_10_,
                         bottom_width_0_height_0_subtile_14__pin_clk_11_,
                         bottom_width_0_height_0_subtile_14__pin_clk_12_,
                         bottom_width_0_height_0_subtile_14__pin_clk_13_,
                         bottom_width_0_height_0_subtile_14__pin_clk_14_,
                         bottom_width_0_height_0_subtile_14__pin_clk_15_,
                         bottom_width_0_height_0_subtile_15__pin_clk_0_,
                         bottom_width_0_height_0_subtile_15__pin_clk_1_,
                         bottom_width_0_height_0_subtile_15__pin_clk_2_,
                         bottom_width_0_height_0_subtile_15__pin_clk_3_,
                         bottom_width_0_height_0_subtile_15__pin_clk_4_,
                         bottom_width_0_height_0_subtile_15__pin_clk_5_,
                         bottom_width_0_height_0_subtile_15__pin_clk_6_,
                         bottom_width_0_height_0_subtile_15__pin_clk_7_,
                         bottom_width_0_height_0_subtile_15__pin_clk_8_,
                         bottom_width_0_height_0_subtile_15__pin_clk_9_,
                         bottom_width_0_height_0_subtile_15__pin_clk_10_,
                         bottom_width_0_height_0_subtile_15__pin_clk_11_,
                         bottom_width_0_height_0_subtile_15__pin_clk_12_,
                         bottom_width_0_height_0_subtile_15__pin_clk_13_,
                         bottom_width_0_height_0_subtile_15__pin_clk_14_,
                         bottom_width_0_height_0_subtile_15__pin_clk_15_,
                         bottom_width_0_height_0_subtile_16__pin_clk_0_,
                         bottom_width_0_height_0_subtile_16__pin_clk_1_,
                         bottom_width_0_height_0_subtile_16__pin_clk_2_,
                         bottom_width_0_height_0_subtile_16__pin_clk_3_,
                         bottom_width_0_height_0_subtile_16__pin_clk_4_,
                         bottom_width_0_height_0_subtile_16__pin_clk_5_,
                         bottom_width_0_height_0_subtile_16__pin_clk_6_,
                         bottom_width_0_height_0_subtile_16__pin_clk_7_,
                         bottom_width_0_height_0_subtile_16__pin_clk_8_,
                         bottom_width_0_height_0_subtile_16__pin_clk_9_,
                         bottom_width_0_height_0_subtile_16__pin_clk_10_,
                         bottom_width_0_height_0_subtile_16__pin_clk_11_,
                         bottom_width_0_height_0_subtile_16__pin_clk_12_,
                         bottom_width_0_height_0_subtile_16__pin_clk_13_,
                         bottom_width_0_height_0_subtile_16__pin_clk_14_,
                         bottom_width_0_height_0_subtile_16__pin_clk_15_,
                         bottom_width_0_height_0_subtile_17__pin_clk_0_,
                         bottom_width_0_height_0_subtile_17__pin_clk_1_,
                         bottom_width_0_height_0_subtile_17__pin_clk_2_,
                         bottom_width_0_height_0_subtile_17__pin_clk_3_,
                         bottom_width_0_height_0_subtile_17__pin_clk_4_,
                         bottom_width_0_height_0_subtile_17__pin_clk_5_,
                         bottom_width_0_height_0_subtile_17__pin_clk_6_,
                         bottom_width_0_height_0_subtile_17__pin_clk_7_,
                         bottom_width_0_height_0_subtile_17__pin_clk_8_,
                         bottom_width_0_height_0_subtile_17__pin_clk_9_,
                         bottom_width_0_height_0_subtile_17__pin_clk_10_,
                         bottom_width_0_height_0_subtile_17__pin_clk_11_,
                         bottom_width_0_height_0_subtile_17__pin_clk_12_,
                         bottom_width_0_height_0_subtile_17__pin_clk_13_,
                         bottom_width_0_height_0_subtile_17__pin_clk_14_,
                         bottom_width_0_height_0_subtile_17__pin_clk_15_,
                         bottom_width_0_height_0_subtile_18__pin_clk_0_,
                         bottom_width_0_height_0_subtile_18__pin_clk_1_,
                         bottom_width_0_height_0_subtile_18__pin_clk_2_,
                         bottom_width_0_height_0_subtile_18__pin_clk_3_,
                         bottom_width_0_height_0_subtile_18__pin_clk_4_,
                         bottom_width_0_height_0_subtile_18__pin_clk_5_,
                         bottom_width_0_height_0_subtile_18__pin_clk_6_,
                         bottom_width_0_height_0_subtile_18__pin_clk_7_,
                         bottom_width_0_height_0_subtile_18__pin_clk_8_,
                         bottom_width_0_height_0_subtile_18__pin_clk_9_,
                         bottom_width_0_height_0_subtile_18__pin_clk_10_,
                         bottom_width_0_height_0_subtile_18__pin_clk_11_,
                         bottom_width_0_height_0_subtile_18__pin_clk_12_,
                         bottom_width_0_height_0_subtile_18__pin_clk_13_,
                         bottom_width_0_height_0_subtile_18__pin_clk_14_,
                         bottom_width_0_height_0_subtile_18__pin_clk_15_,
                         bottom_width_0_height_0_subtile_19__pin_clk_0_,
                         bottom_width_0_height_0_subtile_19__pin_clk_1_,
                         bottom_width_0_height_0_subtile_19__pin_clk_2_,
                         bottom_width_0_height_0_subtile_19__pin_clk_3_,
                         bottom_width_0_height_0_subtile_19__pin_clk_4_,
                         bottom_width_0_height_0_subtile_19__pin_clk_5_,
                         bottom_width_0_height_0_subtile_19__pin_clk_6_,
                         bottom_width_0_height_0_subtile_19__pin_clk_7_,
                         bottom_width_0_height_0_subtile_19__pin_clk_8_,
                         bottom_width_0_height_0_subtile_19__pin_clk_9_,
                         bottom_width_0_height_0_subtile_19__pin_clk_10_,
                         bottom_width_0_height_0_subtile_19__pin_clk_11_,
                         bottom_width_0_height_0_subtile_19__pin_clk_12_,
                         bottom_width_0_height_0_subtile_19__pin_clk_13_,
                         bottom_width_0_height_0_subtile_19__pin_clk_14_,
                         bottom_width_0_height_0_subtile_19__pin_clk_15_,
                         bottom_width_0_height_0_subtile_20__pin_clk_0_,
                         bottom_width_0_height_0_subtile_20__pin_clk_1_,
                         bottom_width_0_height_0_subtile_20__pin_clk_2_,
                         bottom_width_0_height_0_subtile_20__pin_clk_3_,
                         bottom_width_0_height_0_subtile_20__pin_clk_4_,
                         bottom_width_0_height_0_subtile_20__pin_clk_5_,
                         bottom_width_0_height_0_subtile_20__pin_clk_6_,
                         bottom_width_0_height_0_subtile_20__pin_clk_7_,
                         bottom_width_0_height_0_subtile_20__pin_clk_8_,
                         bottom_width_0_height_0_subtile_20__pin_clk_9_,
                         bottom_width_0_height_0_subtile_20__pin_clk_10_,
                         bottom_width_0_height_0_subtile_20__pin_clk_11_,
                         bottom_width_0_height_0_subtile_20__pin_clk_12_,
                         bottom_width_0_height_0_subtile_20__pin_clk_13_,
                         bottom_width_0_height_0_subtile_20__pin_clk_14_,
                         bottom_width_0_height_0_subtile_20__pin_clk_15_,
                         bottom_width_0_height_0_subtile_21__pin_clk_0_,
                         bottom_width_0_height_0_subtile_21__pin_clk_1_,
                         bottom_width_0_height_0_subtile_21__pin_clk_2_,
                         bottom_width_0_height_0_subtile_21__pin_clk_3_,
                         bottom_width_0_height_0_subtile_21__pin_clk_4_,
                         bottom_width_0_height_0_subtile_21__pin_clk_5_,
                         bottom_width_0_height_0_subtile_21__pin_clk_6_,
                         bottom_width_0_height_0_subtile_21__pin_clk_7_,
                         bottom_width_0_height_0_subtile_21__pin_clk_8_,
                         bottom_width_0_height_0_subtile_21__pin_clk_9_,
                         bottom_width_0_height_0_subtile_21__pin_clk_10_,
                         bottom_width_0_height_0_subtile_21__pin_clk_11_,
                         bottom_width_0_height_0_subtile_21__pin_clk_12_,
                         bottom_width_0_height_0_subtile_21__pin_clk_13_,
                         bottom_width_0_height_0_subtile_21__pin_clk_14_,
                         bottom_width_0_height_0_subtile_21__pin_clk_15_,
                         bottom_width_0_height_0_subtile_22__pin_clk_0_,
                         bottom_width_0_height_0_subtile_22__pin_clk_1_,
                         bottom_width_0_height_0_subtile_22__pin_clk_2_,
                         bottom_width_0_height_0_subtile_22__pin_clk_3_,
                         bottom_width_0_height_0_subtile_22__pin_clk_4_,
                         bottom_width_0_height_0_subtile_22__pin_clk_5_,
                         bottom_width_0_height_0_subtile_22__pin_clk_6_,
                         bottom_width_0_height_0_subtile_22__pin_clk_7_,
                         bottom_width_0_height_0_subtile_22__pin_clk_8_,
                         bottom_width_0_height_0_subtile_22__pin_clk_9_,
                         bottom_width_0_height_0_subtile_22__pin_clk_10_,
                         bottom_width_0_height_0_subtile_22__pin_clk_11_,
                         bottom_width_0_height_0_subtile_22__pin_clk_12_,
                         bottom_width_0_height_0_subtile_22__pin_clk_13_,
                         bottom_width_0_height_0_subtile_22__pin_clk_14_,
                         bottom_width_0_height_0_subtile_22__pin_clk_15_,
                         bottom_width_0_height_0_subtile_23__pin_clk_0_,
                         bottom_width_0_height_0_subtile_23__pin_clk_1_,
                         bottom_width_0_height_0_subtile_23__pin_clk_2_,
                         bottom_width_0_height_0_subtile_23__pin_clk_3_,
                         bottom_width_0_height_0_subtile_23__pin_clk_4_,
                         bottom_width_0_height_0_subtile_23__pin_clk_5_,
                         bottom_width_0_height_0_subtile_23__pin_clk_6_,
                         bottom_width_0_height_0_subtile_23__pin_clk_7_,
                         bottom_width_0_height_0_subtile_23__pin_clk_8_,
                         bottom_width_0_height_0_subtile_23__pin_clk_9_,
                         bottom_width_0_height_0_subtile_23__pin_clk_10_,
                         bottom_width_0_height_0_subtile_23__pin_clk_11_,
                         bottom_width_0_height_0_subtile_23__pin_clk_12_,
                         bottom_width_0_height_0_subtile_23__pin_clk_13_,
                         bottom_width_0_height_0_subtile_23__pin_clk_14_,
                         bottom_width_0_height_0_subtile_23__pin_clk_15_,
                         bottom_width_0_height_0_subtile_24__pin_clk_0_,
                         bottom_width_0_height_0_subtile_24__pin_clk_1_,
                         bottom_width_0_height_0_subtile_24__pin_clk_2_,
                         bottom_width_0_height_0_subtile_24__pin_clk_3_,
                         bottom_width_0_height_0_subtile_24__pin_clk_4_,
                         bottom_width_0_height_0_subtile_24__pin_clk_5_,
                         bottom_width_0_height_0_subtile_24__pin_clk_6_,
                         bottom_width_0_height_0_subtile_24__pin_clk_7_,
                         bottom_width_0_height_0_subtile_24__pin_clk_8_,
                         bottom_width_0_height_0_subtile_24__pin_clk_9_,
                         bottom_width_0_height_0_subtile_24__pin_clk_10_,
                         bottom_width_0_height_0_subtile_24__pin_clk_11_,
                         bottom_width_0_height_0_subtile_24__pin_clk_12_,
                         bottom_width_0_height_0_subtile_24__pin_clk_13_,
                         bottom_width_0_height_0_subtile_24__pin_clk_14_,
                         bottom_width_0_height_0_subtile_24__pin_clk_15_,
                         bottom_width_0_height_0_subtile_25__pin_clk_0_,
                         bottom_width_0_height_0_subtile_25__pin_clk_1_,
                         bottom_width_0_height_0_subtile_25__pin_clk_2_,
                         bottom_width_0_height_0_subtile_25__pin_clk_3_,
                         bottom_width_0_height_0_subtile_25__pin_clk_4_,
                         bottom_width_0_height_0_subtile_25__pin_clk_5_,
                         bottom_width_0_height_0_subtile_25__pin_clk_6_,
                         bottom_width_0_height_0_subtile_25__pin_clk_7_,
                         bottom_width_0_height_0_subtile_25__pin_clk_8_,
                         bottom_width_0_height_0_subtile_25__pin_clk_9_,
                         bottom_width_0_height_0_subtile_25__pin_clk_10_,
                         bottom_width_0_height_0_subtile_25__pin_clk_11_,
                         bottom_width_0_height_0_subtile_25__pin_clk_12_,
                         bottom_width_0_height_0_subtile_25__pin_clk_13_,
                         bottom_width_0_height_0_subtile_25__pin_clk_14_,
                         bottom_width_0_height_0_subtile_25__pin_clk_15_,
                         bottom_width_0_height_0_subtile_26__pin_clk_0_,
                         bottom_width_0_height_0_subtile_26__pin_clk_1_,
                         bottom_width_0_height_0_subtile_26__pin_clk_2_,
                         bottom_width_0_height_0_subtile_26__pin_clk_3_,
                         bottom_width_0_height_0_subtile_26__pin_clk_4_,
                         bottom_width_0_height_0_subtile_26__pin_clk_5_,
                         bottom_width_0_height_0_subtile_26__pin_clk_6_,
                         bottom_width_0_height_0_subtile_26__pin_clk_7_,
                         bottom_width_0_height_0_subtile_26__pin_clk_8_,
                         bottom_width_0_height_0_subtile_26__pin_clk_9_,
                         bottom_width_0_height_0_subtile_26__pin_clk_10_,
                         bottom_width_0_height_0_subtile_26__pin_clk_11_,
                         bottom_width_0_height_0_subtile_26__pin_clk_12_,
                         bottom_width_0_height_0_subtile_26__pin_clk_13_,
                         bottom_width_0_height_0_subtile_26__pin_clk_14_,
                         bottom_width_0_height_0_subtile_26__pin_clk_15_,
                         bottom_width_0_height_0_subtile_27__pin_clk_0_,
                         bottom_width_0_height_0_subtile_27__pin_clk_1_,
                         bottom_width_0_height_0_subtile_27__pin_clk_2_,
                         bottom_width_0_height_0_subtile_27__pin_clk_3_,
                         bottom_width_0_height_0_subtile_27__pin_clk_4_,
                         bottom_width_0_height_0_subtile_27__pin_clk_5_,
                         bottom_width_0_height_0_subtile_27__pin_clk_6_,
                         bottom_width_0_height_0_subtile_27__pin_clk_7_,
                         bottom_width_0_height_0_subtile_27__pin_clk_8_,
                         bottom_width_0_height_0_subtile_27__pin_clk_9_,
                         bottom_width_0_height_0_subtile_27__pin_clk_10_,
                         bottom_width_0_height_0_subtile_27__pin_clk_11_,
                         bottom_width_0_height_0_subtile_27__pin_clk_12_,
                         bottom_width_0_height_0_subtile_27__pin_clk_13_,
                         bottom_width_0_height_0_subtile_27__pin_clk_14_,
                         bottom_width_0_height_0_subtile_27__pin_clk_15_,
                         bottom_width_0_height_0_subtile_28__pin_clk_0_,
                         bottom_width_0_height_0_subtile_28__pin_clk_1_,
                         bottom_width_0_height_0_subtile_28__pin_clk_2_,
                         bottom_width_0_height_0_subtile_28__pin_clk_3_,
                         bottom_width_0_height_0_subtile_28__pin_clk_4_,
                         bottom_width_0_height_0_subtile_28__pin_clk_5_,
                         bottom_width_0_height_0_subtile_28__pin_clk_6_,
                         bottom_width_0_height_0_subtile_28__pin_clk_7_,
                         bottom_width_0_height_0_subtile_28__pin_clk_8_,
                         bottom_width_0_height_0_subtile_28__pin_clk_9_,
                         bottom_width_0_height_0_subtile_28__pin_clk_10_,
                         bottom_width_0_height_0_subtile_28__pin_clk_11_,
                         bottom_width_0_height_0_subtile_28__pin_clk_12_,
                         bottom_width_0_height_0_subtile_28__pin_clk_13_,
                         bottom_width_0_height_0_subtile_28__pin_clk_14_,
                         bottom_width_0_height_0_subtile_28__pin_clk_15_,
                         bottom_width_0_height_0_subtile_29__pin_clk_0_,
                         bottom_width_0_height_0_subtile_29__pin_clk_1_,
                         bottom_width_0_height_0_subtile_29__pin_clk_2_,
                         bottom_width_0_height_0_subtile_29__pin_clk_3_,
                         bottom_width_0_height_0_subtile_29__pin_clk_4_,
                         bottom_width_0_height_0_subtile_29__pin_clk_5_,
                         bottom_width_0_height_0_subtile_29__pin_clk_6_,
                         bottom_width_0_height_0_subtile_29__pin_clk_7_,
                         bottom_width_0_height_0_subtile_29__pin_clk_8_,
                         bottom_width_0_height_0_subtile_29__pin_clk_9_,
                         bottom_width_0_height_0_subtile_29__pin_clk_10_,
                         bottom_width_0_height_0_subtile_29__pin_clk_11_,
                         bottom_width_0_height_0_subtile_29__pin_clk_12_,
                         bottom_width_0_height_0_subtile_29__pin_clk_13_,
                         bottom_width_0_height_0_subtile_29__pin_clk_14_,
                         bottom_width_0_height_0_subtile_29__pin_clk_15_,
                         bottom_width_0_height_0_subtile_30__pin_clk_0_,
                         bottom_width_0_height_0_subtile_30__pin_clk_1_,
                         bottom_width_0_height_0_subtile_30__pin_clk_2_,
                         bottom_width_0_height_0_subtile_30__pin_clk_3_,
                         bottom_width_0_height_0_subtile_30__pin_clk_4_,
                         bottom_width_0_height_0_subtile_30__pin_clk_5_,
                         bottom_width_0_height_0_subtile_30__pin_clk_6_,
                         bottom_width_0_height_0_subtile_30__pin_clk_7_,
                         bottom_width_0_height_0_subtile_30__pin_clk_8_,
                         bottom_width_0_height_0_subtile_30__pin_clk_9_,
                         bottom_width_0_height_0_subtile_30__pin_clk_10_,
                         bottom_width_0_height_0_subtile_30__pin_clk_11_,
                         bottom_width_0_height_0_subtile_30__pin_clk_12_,
                         bottom_width_0_height_0_subtile_30__pin_clk_13_,
                         bottom_width_0_height_0_subtile_30__pin_clk_14_,
                         bottom_width_0_height_0_subtile_30__pin_clk_15_,
                         bottom_width_0_height_0_subtile_31__pin_clk_0_,
                         bottom_width_0_height_0_subtile_31__pin_clk_1_,
                         bottom_width_0_height_0_subtile_31__pin_clk_2_,
                         bottom_width_0_height_0_subtile_31__pin_clk_3_,
                         bottom_width_0_height_0_subtile_31__pin_clk_4_,
                         bottom_width_0_height_0_subtile_31__pin_clk_5_,
                         bottom_width_0_height_0_subtile_31__pin_clk_6_,
                         bottom_width_0_height_0_subtile_31__pin_clk_7_,
                         bottom_width_0_height_0_subtile_31__pin_clk_8_,
                         bottom_width_0_height_0_subtile_31__pin_clk_9_,
                         bottom_width_0_height_0_subtile_31__pin_clk_10_,
                         bottom_width_0_height_0_subtile_31__pin_clk_11_,
                         bottom_width_0_height_0_subtile_31__pin_clk_12_,
                         bottom_width_0_height_0_subtile_31__pin_clk_13_,
                         bottom_width_0_height_0_subtile_31__pin_clk_14_,
                         bottom_width_0_height_0_subtile_31__pin_clk_15_,
                         bottom_width_0_height_0_subtile_32__pin_clk_0_,
                         bottom_width_0_height_0_subtile_32__pin_clk_1_,
                         bottom_width_0_height_0_subtile_32__pin_clk_2_,
                         bottom_width_0_height_0_subtile_32__pin_clk_3_,
                         bottom_width_0_height_0_subtile_32__pin_clk_4_,
                         bottom_width_0_height_0_subtile_32__pin_clk_5_,
                         bottom_width_0_height_0_subtile_32__pin_clk_6_,
                         bottom_width_0_height_0_subtile_32__pin_clk_7_,
                         bottom_width_0_height_0_subtile_32__pin_clk_8_,
                         bottom_width_0_height_0_subtile_32__pin_clk_9_,
                         bottom_width_0_height_0_subtile_32__pin_clk_10_,
                         bottom_width_0_height_0_subtile_32__pin_clk_11_,
                         bottom_width_0_height_0_subtile_32__pin_clk_12_,
                         bottom_width_0_height_0_subtile_32__pin_clk_13_,
                         bottom_width_0_height_0_subtile_32__pin_clk_14_,
                         bottom_width_0_height_0_subtile_32__pin_clk_15_,
                         bottom_width_0_height_0_subtile_33__pin_clk_0_,
                         bottom_width_0_height_0_subtile_33__pin_clk_1_,
                         bottom_width_0_height_0_subtile_33__pin_clk_2_,
                         bottom_width_0_height_0_subtile_33__pin_clk_3_,
                         bottom_width_0_height_0_subtile_33__pin_clk_4_,
                         bottom_width_0_height_0_subtile_33__pin_clk_5_,
                         bottom_width_0_height_0_subtile_33__pin_clk_6_,
                         bottom_width_0_height_0_subtile_33__pin_clk_7_,
                         bottom_width_0_height_0_subtile_33__pin_clk_8_,
                         bottom_width_0_height_0_subtile_33__pin_clk_9_,
                         bottom_width_0_height_0_subtile_33__pin_clk_10_,
                         bottom_width_0_height_0_subtile_33__pin_clk_11_,
                         bottom_width_0_height_0_subtile_33__pin_clk_12_,
                         bottom_width_0_height_0_subtile_33__pin_clk_13_,
                         bottom_width_0_height_0_subtile_33__pin_clk_14_,
                         bottom_width_0_height_0_subtile_33__pin_clk_15_,
                         bottom_width_0_height_0_subtile_34__pin_clk_0_,
                         bottom_width_0_height_0_subtile_34__pin_clk_1_,
                         bottom_width_0_height_0_subtile_34__pin_clk_2_,
                         bottom_width_0_height_0_subtile_34__pin_clk_3_,
                         bottom_width_0_height_0_subtile_34__pin_clk_4_,
                         bottom_width_0_height_0_subtile_34__pin_clk_5_,
                         bottom_width_0_height_0_subtile_34__pin_clk_6_,
                         bottom_width_0_height_0_subtile_34__pin_clk_7_,
                         bottom_width_0_height_0_subtile_34__pin_clk_8_,
                         bottom_width_0_height_0_subtile_34__pin_clk_9_,
                         bottom_width_0_height_0_subtile_34__pin_clk_10_,
                         bottom_width_0_height_0_subtile_34__pin_clk_11_,
                         bottom_width_0_height_0_subtile_34__pin_clk_12_,
                         bottom_width_0_height_0_subtile_34__pin_clk_13_,
                         bottom_width_0_height_0_subtile_34__pin_clk_14_,
                         bottom_width_0_height_0_subtile_34__pin_clk_15_,
                         bottom_width_0_height_0_subtile_35__pin_clk_0_,
                         bottom_width_0_height_0_subtile_35__pin_clk_1_,
                         bottom_width_0_height_0_subtile_35__pin_clk_2_,
                         bottom_width_0_height_0_subtile_35__pin_clk_3_,
                         bottom_width_0_height_0_subtile_35__pin_clk_4_,
                         bottom_width_0_height_0_subtile_35__pin_clk_5_,
                         bottom_width_0_height_0_subtile_35__pin_clk_6_,
                         bottom_width_0_height_0_subtile_35__pin_clk_7_,
                         bottom_width_0_height_0_subtile_35__pin_clk_8_,
                         bottom_width_0_height_0_subtile_35__pin_clk_9_,
                         bottom_width_0_height_0_subtile_35__pin_clk_10_,
                         bottom_width_0_height_0_subtile_35__pin_clk_11_,
                         bottom_width_0_height_0_subtile_35__pin_clk_12_,
                         bottom_width_0_height_0_subtile_35__pin_clk_13_,
                         bottom_width_0_height_0_subtile_35__pin_clk_14_,
                         bottom_width_0_height_0_subtile_35__pin_clk_15_,
                         bottom_width_0_height_0_subtile_36__pin_clk_0_,
                         bottom_width_0_height_0_subtile_36__pin_clk_1_,
                         bottom_width_0_height_0_subtile_36__pin_clk_2_,
                         bottom_width_0_height_0_subtile_36__pin_clk_3_,
                         bottom_width_0_height_0_subtile_36__pin_clk_4_,
                         bottom_width_0_height_0_subtile_36__pin_clk_5_,
                         bottom_width_0_height_0_subtile_36__pin_clk_6_,
                         bottom_width_0_height_0_subtile_36__pin_clk_7_,
                         bottom_width_0_height_0_subtile_36__pin_clk_8_,
                         bottom_width_0_height_0_subtile_36__pin_clk_9_,
                         bottom_width_0_height_0_subtile_36__pin_clk_10_,
                         bottom_width_0_height_0_subtile_36__pin_clk_11_,
                         bottom_width_0_height_0_subtile_36__pin_clk_12_,
                         bottom_width_0_height_0_subtile_36__pin_clk_13_,
                         bottom_width_0_height_0_subtile_36__pin_clk_14_,
                         bottom_width_0_height_0_subtile_36__pin_clk_15_,
                         bottom_width_0_height_0_subtile_37__pin_clk_0_,
                         bottom_width_0_height_0_subtile_37__pin_clk_1_,
                         bottom_width_0_height_0_subtile_37__pin_clk_2_,
                         bottom_width_0_height_0_subtile_37__pin_clk_3_,
                         bottom_width_0_height_0_subtile_37__pin_clk_4_,
                         bottom_width_0_height_0_subtile_37__pin_clk_5_,
                         bottom_width_0_height_0_subtile_37__pin_clk_6_,
                         bottom_width_0_height_0_subtile_37__pin_clk_7_,
                         bottom_width_0_height_0_subtile_37__pin_clk_8_,
                         bottom_width_0_height_0_subtile_37__pin_clk_9_,
                         bottom_width_0_height_0_subtile_37__pin_clk_10_,
                         bottom_width_0_height_0_subtile_37__pin_clk_11_,
                         bottom_width_0_height_0_subtile_37__pin_clk_12_,
                         bottom_width_0_height_0_subtile_37__pin_clk_13_,
                         bottom_width_0_height_0_subtile_37__pin_clk_14_,
                         bottom_width_0_height_0_subtile_37__pin_clk_15_,
                         bottom_width_0_height_0_subtile_38__pin_clk_0_,
                         bottom_width_0_height_0_subtile_38__pin_clk_1_,
                         bottom_width_0_height_0_subtile_38__pin_clk_2_,
                         bottom_width_0_height_0_subtile_38__pin_clk_3_,
                         bottom_width_0_height_0_subtile_38__pin_clk_4_,
                         bottom_width_0_height_0_subtile_38__pin_clk_5_,
                         bottom_width_0_height_0_subtile_38__pin_clk_6_,
                         bottom_width_0_height_0_subtile_38__pin_clk_7_,
                         bottom_width_0_height_0_subtile_38__pin_clk_8_,
                         bottom_width_0_height_0_subtile_38__pin_clk_9_,
                         bottom_width_0_height_0_subtile_38__pin_clk_10_,
                         bottom_width_0_height_0_subtile_38__pin_clk_11_,
                         bottom_width_0_height_0_subtile_38__pin_clk_12_,
                         bottom_width_0_height_0_subtile_38__pin_clk_13_,
                         bottom_width_0_height_0_subtile_38__pin_clk_14_,
                         bottom_width_0_height_0_subtile_38__pin_clk_15_,
                         bottom_width_0_height_0_subtile_39__pin_clk_0_,
                         bottom_width_0_height_0_subtile_39__pin_clk_1_,
                         bottom_width_0_height_0_subtile_39__pin_clk_2_,
                         bottom_width_0_height_0_subtile_39__pin_clk_3_,
                         bottom_width_0_height_0_subtile_39__pin_clk_4_,
                         bottom_width_0_height_0_subtile_39__pin_clk_5_,
                         bottom_width_0_height_0_subtile_39__pin_clk_6_,
                         bottom_width_0_height_0_subtile_39__pin_clk_7_,
                         bottom_width_0_height_0_subtile_39__pin_clk_8_,
                         bottom_width_0_height_0_subtile_39__pin_clk_9_,
                         bottom_width_0_height_0_subtile_39__pin_clk_10_,
                         bottom_width_0_height_0_subtile_39__pin_clk_11_,
                         bottom_width_0_height_0_subtile_39__pin_clk_12_,
                         bottom_width_0_height_0_subtile_39__pin_clk_13_,
                         bottom_width_0_height_0_subtile_39__pin_clk_14_,
                         bottom_width_0_height_0_subtile_39__pin_clk_15_,
                         bottom_width_0_height_0_subtile_40__pin_clk_0_,
                         bottom_width_0_height_0_subtile_40__pin_clk_1_,
                         bottom_width_0_height_0_subtile_40__pin_clk_2_,
                         bottom_width_0_height_0_subtile_40__pin_clk_3_,
                         bottom_width_0_height_0_subtile_40__pin_clk_4_,
                         bottom_width_0_height_0_subtile_40__pin_clk_5_,
                         bottom_width_0_height_0_subtile_40__pin_clk_6_,
                         bottom_width_0_height_0_subtile_40__pin_clk_7_,
                         bottom_width_0_height_0_subtile_40__pin_clk_8_,
                         bottom_width_0_height_0_subtile_40__pin_clk_9_,
                         bottom_width_0_height_0_subtile_40__pin_clk_10_,
                         bottom_width_0_height_0_subtile_40__pin_clk_11_,
                         bottom_width_0_height_0_subtile_40__pin_clk_12_,
                         bottom_width_0_height_0_subtile_40__pin_clk_13_,
                         bottom_width_0_height_0_subtile_40__pin_clk_14_,
                         bottom_width_0_height_0_subtile_40__pin_clk_15_,
                         bottom_width_0_height_0_subtile_41__pin_clk_0_,
                         bottom_width_0_height_0_subtile_41__pin_clk_1_,
                         bottom_width_0_height_0_subtile_41__pin_clk_2_,
                         bottom_width_0_height_0_subtile_41__pin_clk_3_,
                         bottom_width_0_height_0_subtile_41__pin_clk_4_,
                         bottom_width_0_height_0_subtile_41__pin_clk_5_,
                         bottom_width_0_height_0_subtile_41__pin_clk_6_,
                         bottom_width_0_height_0_subtile_41__pin_clk_7_,
                         bottom_width_0_height_0_subtile_41__pin_clk_8_,
                         bottom_width_0_height_0_subtile_41__pin_clk_9_,
                         bottom_width_0_height_0_subtile_41__pin_clk_10_,
                         bottom_width_0_height_0_subtile_41__pin_clk_11_,
                         bottom_width_0_height_0_subtile_41__pin_clk_12_,
                         bottom_width_0_height_0_subtile_41__pin_clk_13_,
                         bottom_width_0_height_0_subtile_41__pin_clk_14_,
                         bottom_width_0_height_0_subtile_41__pin_clk_15_,
                         bottom_width_0_height_0_subtile_42__pin_clk_0_,
                         bottom_width_0_height_0_subtile_42__pin_clk_1_,
                         bottom_width_0_height_0_subtile_42__pin_clk_2_,
                         bottom_width_0_height_0_subtile_42__pin_clk_3_,
                         bottom_width_0_height_0_subtile_42__pin_clk_4_,
                         bottom_width_0_height_0_subtile_42__pin_clk_5_,
                         bottom_width_0_height_0_subtile_42__pin_clk_6_,
                         bottom_width_0_height_0_subtile_42__pin_clk_7_,
                         bottom_width_0_height_0_subtile_42__pin_clk_8_,
                         bottom_width_0_height_0_subtile_42__pin_clk_9_,
                         bottom_width_0_height_0_subtile_42__pin_clk_10_,
                         bottom_width_0_height_0_subtile_42__pin_clk_11_,
                         bottom_width_0_height_0_subtile_42__pin_clk_12_,
                         bottom_width_0_height_0_subtile_42__pin_clk_13_,
                         bottom_width_0_height_0_subtile_42__pin_clk_14_,
                         bottom_width_0_height_0_subtile_42__pin_clk_15_,
                         bottom_width_0_height_0_subtile_43__pin_clk_0_,
                         bottom_width_0_height_0_subtile_43__pin_clk_1_,
                         bottom_width_0_height_0_subtile_43__pin_clk_2_,
                         bottom_width_0_height_0_subtile_43__pin_clk_3_,
                         bottom_width_0_height_0_subtile_43__pin_clk_4_,
                         bottom_width_0_height_0_subtile_43__pin_clk_5_,
                         bottom_width_0_height_0_subtile_43__pin_clk_6_,
                         bottom_width_0_height_0_subtile_43__pin_clk_7_,
                         bottom_width_0_height_0_subtile_43__pin_clk_8_,
                         bottom_width_0_height_0_subtile_43__pin_clk_9_,
                         bottom_width_0_height_0_subtile_43__pin_clk_10_,
                         bottom_width_0_height_0_subtile_43__pin_clk_11_,
                         bottom_width_0_height_0_subtile_43__pin_clk_12_,
                         bottom_width_0_height_0_subtile_43__pin_clk_13_,
                         bottom_width_0_height_0_subtile_43__pin_clk_14_,
                         bottom_width_0_height_0_subtile_43__pin_clk_15_,
                         bottom_width_0_height_0_subtile_44__pin_clk_0_,
                         bottom_width_0_height_0_subtile_44__pin_clk_1_,
                         bottom_width_0_height_0_subtile_44__pin_clk_2_,
                         bottom_width_0_height_0_subtile_44__pin_clk_3_,
                         bottom_width_0_height_0_subtile_44__pin_clk_4_,
                         bottom_width_0_height_0_subtile_44__pin_clk_5_,
                         bottom_width_0_height_0_subtile_44__pin_clk_6_,
                         bottom_width_0_height_0_subtile_44__pin_clk_7_,
                         bottom_width_0_height_0_subtile_44__pin_clk_8_,
                         bottom_width_0_height_0_subtile_44__pin_clk_9_,
                         bottom_width_0_height_0_subtile_44__pin_clk_10_,
                         bottom_width_0_height_0_subtile_44__pin_clk_11_,
                         bottom_width_0_height_0_subtile_44__pin_clk_12_,
                         bottom_width_0_height_0_subtile_44__pin_clk_13_,
                         bottom_width_0_height_0_subtile_44__pin_clk_14_,
                         bottom_width_0_height_0_subtile_44__pin_clk_15_,
                         bottom_width_0_height_0_subtile_45__pin_clk_0_,
                         bottom_width_0_height_0_subtile_45__pin_clk_1_,
                         bottom_width_0_height_0_subtile_45__pin_clk_2_,
                         bottom_width_0_height_0_subtile_45__pin_clk_3_,
                         bottom_width_0_height_0_subtile_45__pin_clk_4_,
                         bottom_width_0_height_0_subtile_45__pin_clk_5_,
                         bottom_width_0_height_0_subtile_45__pin_clk_6_,
                         bottom_width_0_height_0_subtile_45__pin_clk_7_,
                         bottom_width_0_height_0_subtile_45__pin_clk_8_,
                         bottom_width_0_height_0_subtile_45__pin_clk_9_,
                         bottom_width_0_height_0_subtile_45__pin_clk_10_,
                         bottom_width_0_height_0_subtile_45__pin_clk_11_,
                         bottom_width_0_height_0_subtile_45__pin_clk_12_,
                         bottom_width_0_height_0_subtile_45__pin_clk_13_,
                         bottom_width_0_height_0_subtile_45__pin_clk_14_,
                         bottom_width_0_height_0_subtile_45__pin_clk_15_,
                         bottom_width_0_height_0_subtile_46__pin_clk_0_,
                         bottom_width_0_height_0_subtile_46__pin_clk_1_,
                         bottom_width_0_height_0_subtile_46__pin_clk_2_,
                         bottom_width_0_height_0_subtile_46__pin_clk_3_,
                         bottom_width_0_height_0_subtile_46__pin_clk_4_,
                         bottom_width_0_height_0_subtile_46__pin_clk_5_,
                         bottom_width_0_height_0_subtile_46__pin_clk_6_,
                         bottom_width_0_height_0_subtile_46__pin_clk_7_,
                         bottom_width_0_height_0_subtile_46__pin_clk_8_,
                         bottom_width_0_height_0_subtile_46__pin_clk_9_,
                         bottom_width_0_height_0_subtile_46__pin_clk_10_,
                         bottom_width_0_height_0_subtile_46__pin_clk_11_,
                         bottom_width_0_height_0_subtile_46__pin_clk_12_,
                         bottom_width_0_height_0_subtile_46__pin_clk_13_,
                         bottom_width_0_height_0_subtile_46__pin_clk_14_,
                         bottom_width_0_height_0_subtile_46__pin_clk_15_,
                         bottom_width_0_height_0_subtile_47__pin_clk_0_,
                         bottom_width_0_height_0_subtile_47__pin_clk_1_,
                         bottom_width_0_height_0_subtile_47__pin_clk_2_,
                         bottom_width_0_height_0_subtile_47__pin_clk_3_,
                         bottom_width_0_height_0_subtile_47__pin_clk_4_,
                         bottom_width_0_height_0_subtile_47__pin_clk_5_,
                         bottom_width_0_height_0_subtile_47__pin_clk_6_,
                         bottom_width_0_height_0_subtile_47__pin_clk_7_,
                         bottom_width_0_height_0_subtile_47__pin_clk_8_,
                         bottom_width_0_height_0_subtile_47__pin_clk_9_,
                         bottom_width_0_height_0_subtile_47__pin_clk_10_,
                         bottom_width_0_height_0_subtile_47__pin_clk_11_,
                         bottom_width_0_height_0_subtile_47__pin_clk_12_,
                         bottom_width_0_height_0_subtile_47__pin_clk_13_,
                         bottom_width_0_height_0_subtile_47__pin_clk_14_,
                         bottom_width_0_height_0_subtile_47__pin_clk_15_,
                         bottom_width_0_height_0_subtile_48__pin_clk_0_,
                         bottom_width_0_height_0_subtile_48__pin_clk_1_,
                         bottom_width_0_height_0_subtile_48__pin_clk_2_,
                         bottom_width_0_height_0_subtile_48__pin_clk_3_,
                         bottom_width_0_height_0_subtile_48__pin_clk_4_,
                         bottom_width_0_height_0_subtile_48__pin_clk_5_,
                         bottom_width_0_height_0_subtile_48__pin_clk_6_,
                         bottom_width_0_height_0_subtile_48__pin_clk_7_,
                         bottom_width_0_height_0_subtile_48__pin_clk_8_,
                         bottom_width_0_height_0_subtile_48__pin_clk_9_,
                         bottom_width_0_height_0_subtile_48__pin_clk_10_,
                         bottom_width_0_height_0_subtile_48__pin_clk_11_,
                         bottom_width_0_height_0_subtile_48__pin_clk_12_,
                         bottom_width_0_height_0_subtile_48__pin_clk_13_,
                         bottom_width_0_height_0_subtile_48__pin_clk_14_,
                         bottom_width_0_height_0_subtile_48__pin_clk_15_,
                         bottom_width_0_height_0_subtile_49__pin_clk_0_,
                         bottom_width_0_height_0_subtile_49__pin_clk_1_,
                         bottom_width_0_height_0_subtile_49__pin_clk_2_,
                         bottom_width_0_height_0_subtile_49__pin_clk_3_,
                         bottom_width_0_height_0_subtile_49__pin_clk_4_,
                         bottom_width_0_height_0_subtile_49__pin_clk_5_,
                         bottom_width_0_height_0_subtile_49__pin_clk_6_,
                         bottom_width_0_height_0_subtile_49__pin_clk_7_,
                         bottom_width_0_height_0_subtile_49__pin_clk_8_,
                         bottom_width_0_height_0_subtile_49__pin_clk_9_,
                         bottom_width_0_height_0_subtile_49__pin_clk_10_,
                         bottom_width_0_height_0_subtile_49__pin_clk_11_,
                         bottom_width_0_height_0_subtile_49__pin_clk_12_,
                         bottom_width_0_height_0_subtile_49__pin_clk_13_,
                         bottom_width_0_height_0_subtile_49__pin_clk_14_,
                         bottom_width_0_height_0_subtile_49__pin_clk_15_,
                         bottom_width_0_height_0_subtile_50__pin_clk_0_,
                         bottom_width_0_height_0_subtile_50__pin_clk_1_,
                         bottom_width_0_height_0_subtile_50__pin_clk_2_,
                         bottom_width_0_height_0_subtile_50__pin_clk_3_,
                         bottom_width_0_height_0_subtile_50__pin_clk_4_,
                         bottom_width_0_height_0_subtile_50__pin_clk_5_,
                         bottom_width_0_height_0_subtile_50__pin_clk_6_,
                         bottom_width_0_height_0_subtile_50__pin_clk_7_,
                         bottom_width_0_height_0_subtile_50__pin_clk_8_,
                         bottom_width_0_height_0_subtile_50__pin_clk_9_,
                         bottom_width_0_height_0_subtile_50__pin_clk_10_,
                         bottom_width_0_height_0_subtile_50__pin_clk_11_,
                         bottom_width_0_height_0_subtile_50__pin_clk_12_,
                         bottom_width_0_height_0_subtile_50__pin_clk_13_,
                         bottom_width_0_height_0_subtile_50__pin_clk_14_,
                         bottom_width_0_height_0_subtile_50__pin_clk_15_,
                         bottom_width_0_height_0_subtile_51__pin_clk_0_,
                         bottom_width_0_height_0_subtile_51__pin_clk_1_,
                         bottom_width_0_height_0_subtile_51__pin_clk_2_,
                         bottom_width_0_height_0_subtile_51__pin_clk_3_,
                         bottom_width_0_height_0_subtile_51__pin_clk_4_,
                         bottom_width_0_height_0_subtile_51__pin_clk_5_,
                         bottom_width_0_height_0_subtile_51__pin_clk_6_,
                         bottom_width_0_height_0_subtile_51__pin_clk_7_,
                         bottom_width_0_height_0_subtile_51__pin_clk_8_,
                         bottom_width_0_height_0_subtile_51__pin_clk_9_,
                         bottom_width_0_height_0_subtile_51__pin_clk_10_,
                         bottom_width_0_height_0_subtile_51__pin_clk_11_,
                         bottom_width_0_height_0_subtile_51__pin_clk_12_,
                         bottom_width_0_height_0_subtile_51__pin_clk_13_,
                         bottom_width_0_height_0_subtile_51__pin_clk_14_,
                         bottom_width_0_height_0_subtile_51__pin_clk_15_,
                         bottom_width_0_height_0_subtile_52__pin_clk_0_,
                         bottom_width_0_height_0_subtile_52__pin_clk_1_,
                         bottom_width_0_height_0_subtile_52__pin_clk_2_,
                         bottom_width_0_height_0_subtile_52__pin_clk_3_,
                         bottom_width_0_height_0_subtile_52__pin_clk_4_,
                         bottom_width_0_height_0_subtile_52__pin_clk_5_,
                         bottom_width_0_height_0_subtile_52__pin_clk_6_,
                         bottom_width_0_height_0_subtile_52__pin_clk_7_,
                         bottom_width_0_height_0_subtile_52__pin_clk_8_,
                         bottom_width_0_height_0_subtile_52__pin_clk_9_,
                         bottom_width_0_height_0_subtile_52__pin_clk_10_,
                         bottom_width_0_height_0_subtile_52__pin_clk_11_,
                         bottom_width_0_height_0_subtile_52__pin_clk_12_,
                         bottom_width_0_height_0_subtile_52__pin_clk_13_,
                         bottom_width_0_height_0_subtile_52__pin_clk_14_,
                         bottom_width_0_height_0_subtile_52__pin_clk_15_,
                         bottom_width_0_height_0_subtile_53__pin_clk_0_,
                         bottom_width_0_height_0_subtile_53__pin_clk_1_,
                         bottom_width_0_height_0_subtile_53__pin_clk_2_,
                         bottom_width_0_height_0_subtile_53__pin_clk_3_,
                         bottom_width_0_height_0_subtile_53__pin_clk_4_,
                         bottom_width_0_height_0_subtile_53__pin_clk_5_,
                         bottom_width_0_height_0_subtile_53__pin_clk_6_,
                         bottom_width_0_height_0_subtile_53__pin_clk_7_,
                         bottom_width_0_height_0_subtile_53__pin_clk_8_,
                         bottom_width_0_height_0_subtile_53__pin_clk_9_,
                         bottom_width_0_height_0_subtile_53__pin_clk_10_,
                         bottom_width_0_height_0_subtile_53__pin_clk_11_,
                         bottom_width_0_height_0_subtile_53__pin_clk_12_,
                         bottom_width_0_height_0_subtile_53__pin_clk_13_,
                         bottom_width_0_height_0_subtile_53__pin_clk_14_,
                         bottom_width_0_height_0_subtile_53__pin_clk_15_,
                         bottom_width_0_height_0_subtile_54__pin_clk_0_,
                         bottom_width_0_height_0_subtile_54__pin_clk_1_,
                         bottom_width_0_height_0_subtile_54__pin_clk_2_,
                         bottom_width_0_height_0_subtile_54__pin_clk_3_,
                         bottom_width_0_height_0_subtile_54__pin_clk_4_,
                         bottom_width_0_height_0_subtile_54__pin_clk_5_,
                         bottom_width_0_height_0_subtile_54__pin_clk_6_,
                         bottom_width_0_height_0_subtile_54__pin_clk_7_,
                         bottom_width_0_height_0_subtile_54__pin_clk_8_,
                         bottom_width_0_height_0_subtile_54__pin_clk_9_,
                         bottom_width_0_height_0_subtile_54__pin_clk_10_,
                         bottom_width_0_height_0_subtile_54__pin_clk_11_,
                         bottom_width_0_height_0_subtile_54__pin_clk_12_,
                         bottom_width_0_height_0_subtile_54__pin_clk_13_,
                         bottom_width_0_height_0_subtile_54__pin_clk_14_,
                         bottom_width_0_height_0_subtile_54__pin_clk_15_,
                         bottom_width_0_height_0_subtile_55__pin_clk_0_,
                         bottom_width_0_height_0_subtile_55__pin_clk_1_,
                         bottom_width_0_height_0_subtile_55__pin_clk_2_,
                         bottom_width_0_height_0_subtile_55__pin_clk_3_,
                         bottom_width_0_height_0_subtile_55__pin_clk_4_,
                         bottom_width_0_height_0_subtile_55__pin_clk_5_,
                         bottom_width_0_height_0_subtile_55__pin_clk_6_,
                         bottom_width_0_height_0_subtile_55__pin_clk_7_,
                         bottom_width_0_height_0_subtile_55__pin_clk_8_,
                         bottom_width_0_height_0_subtile_55__pin_clk_9_,
                         bottom_width_0_height_0_subtile_55__pin_clk_10_,
                         bottom_width_0_height_0_subtile_55__pin_clk_11_,
                         bottom_width_0_height_0_subtile_55__pin_clk_12_,
                         bottom_width_0_height_0_subtile_55__pin_clk_13_,
                         bottom_width_0_height_0_subtile_55__pin_clk_14_,
                         bottom_width_0_height_0_subtile_55__pin_clk_15_,
                         bottom_width_0_height_0_subtile_56__pin_clk_0_,
                         bottom_width_0_height_0_subtile_56__pin_clk_1_,
                         bottom_width_0_height_0_subtile_56__pin_clk_2_,
                         bottom_width_0_height_0_subtile_56__pin_clk_3_,
                         bottom_width_0_height_0_subtile_56__pin_clk_4_,
                         bottom_width_0_height_0_subtile_56__pin_clk_5_,
                         bottom_width_0_height_0_subtile_56__pin_clk_6_,
                         bottom_width_0_height_0_subtile_56__pin_clk_7_,
                         bottom_width_0_height_0_subtile_56__pin_clk_8_,
                         bottom_width_0_height_0_subtile_56__pin_clk_9_,
                         bottom_width_0_height_0_subtile_56__pin_clk_10_,
                         bottom_width_0_height_0_subtile_56__pin_clk_11_,
                         bottom_width_0_height_0_subtile_56__pin_clk_12_,
                         bottom_width_0_height_0_subtile_56__pin_clk_13_,
                         bottom_width_0_height_0_subtile_56__pin_clk_14_,
                         bottom_width_0_height_0_subtile_56__pin_clk_15_,
                         bottom_width_0_height_0_subtile_57__pin_clk_0_,
                         bottom_width_0_height_0_subtile_57__pin_clk_1_,
                         bottom_width_0_height_0_subtile_57__pin_clk_2_,
                         bottom_width_0_height_0_subtile_57__pin_clk_3_,
                         bottom_width_0_height_0_subtile_57__pin_clk_4_,
                         bottom_width_0_height_0_subtile_57__pin_clk_5_,
                         bottom_width_0_height_0_subtile_57__pin_clk_6_,
                         bottom_width_0_height_0_subtile_57__pin_clk_7_,
                         bottom_width_0_height_0_subtile_57__pin_clk_8_,
                         bottom_width_0_height_0_subtile_57__pin_clk_9_,
                         bottom_width_0_height_0_subtile_57__pin_clk_10_,
                         bottom_width_0_height_0_subtile_57__pin_clk_11_,
                         bottom_width_0_height_0_subtile_57__pin_clk_12_,
                         bottom_width_0_height_0_subtile_57__pin_clk_13_,
                         bottom_width_0_height_0_subtile_57__pin_clk_14_,
                         bottom_width_0_height_0_subtile_57__pin_clk_15_,
                         bottom_width_0_height_0_subtile_58__pin_clk_0_,
                         bottom_width_0_height_0_subtile_58__pin_clk_1_,
                         bottom_width_0_height_0_subtile_58__pin_clk_2_,
                         bottom_width_0_height_0_subtile_58__pin_clk_3_,
                         bottom_width_0_height_0_subtile_58__pin_clk_4_,
                         bottom_width_0_height_0_subtile_58__pin_clk_5_,
                         bottom_width_0_height_0_subtile_58__pin_clk_6_,
                         bottom_width_0_height_0_subtile_58__pin_clk_7_,
                         bottom_width_0_height_0_subtile_58__pin_clk_8_,
                         bottom_width_0_height_0_subtile_58__pin_clk_9_,
                         bottom_width_0_height_0_subtile_58__pin_clk_10_,
                         bottom_width_0_height_0_subtile_58__pin_clk_11_,
                         bottom_width_0_height_0_subtile_58__pin_clk_12_,
                         bottom_width_0_height_0_subtile_58__pin_clk_13_,
                         bottom_width_0_height_0_subtile_58__pin_clk_14_,
                         bottom_width_0_height_0_subtile_58__pin_clk_15_,
                         bottom_width_0_height_0_subtile_59__pin_clk_0_,
                         bottom_width_0_height_0_subtile_59__pin_clk_1_,
                         bottom_width_0_height_0_subtile_59__pin_clk_2_,
                         bottom_width_0_height_0_subtile_59__pin_clk_3_,
                         bottom_width_0_height_0_subtile_59__pin_clk_4_,
                         bottom_width_0_height_0_subtile_59__pin_clk_5_,
                         bottom_width_0_height_0_subtile_59__pin_clk_6_,
                         bottom_width_0_height_0_subtile_59__pin_clk_7_,
                         bottom_width_0_height_0_subtile_59__pin_clk_8_,
                         bottom_width_0_height_0_subtile_59__pin_clk_9_,
                         bottom_width_0_height_0_subtile_59__pin_clk_10_,
                         bottom_width_0_height_0_subtile_59__pin_clk_11_,
                         bottom_width_0_height_0_subtile_59__pin_clk_12_,
                         bottom_width_0_height_0_subtile_59__pin_clk_13_,
                         bottom_width_0_height_0_subtile_59__pin_clk_14_,
                         bottom_width_0_height_0_subtile_59__pin_clk_15_,
                         left_width_0_height_0_subtile_0__pin_sc_in_0_,
                         left_width_0_height_0_subtile_1__pin_sc_in_0_,
                         left_width_0_height_0_subtile_2__pin_sc_in_0_,
                         left_width_0_height_0_subtile_3__pin_sc_in_0_,
                         left_width_0_height_0_subtile_4__pin_sc_in_0_,
                         left_width_0_height_0_subtile_5__pin_sc_in_0_,
                         left_width_0_height_0_subtile_6__pin_sc_in_0_,
                         left_width_0_height_0_subtile_7__pin_sc_in_0_,
                         left_width_0_height_0_subtile_8__pin_sc_in_0_,
                         left_width_0_height_0_subtile_9__pin_sc_in_0_,
                         left_width_0_height_0_subtile_10__pin_sc_in_0_,
                         left_width_0_height_0_subtile_11__pin_sc_in_0_,
                         left_width_0_height_0_subtile_12__pin_sc_in_0_,
                         left_width_0_height_0_subtile_13__pin_sc_in_0_,
                         left_width_0_height_0_subtile_14__pin_sc_in_0_,
                         left_width_0_height_0_subtile_15__pin_sc_in_0_,
                         left_width_0_height_0_subtile_16__pin_sc_in_0_,
                         left_width_0_height_0_subtile_17__pin_sc_in_0_,
                         left_width_0_height_0_subtile_18__pin_sc_in_0_,
                         left_width_0_height_0_subtile_19__pin_sc_in_0_,
                         left_width_0_height_0_subtile_20__pin_sc_in_0_,
                         left_width_0_height_0_subtile_21__pin_sc_in_0_,
                         left_width_0_height_0_subtile_22__pin_sc_in_0_,
                         left_width_0_height_0_subtile_23__pin_sc_in_0_,
                         left_width_0_height_0_subtile_24__pin_sc_in_0_,
                         left_width_0_height_0_subtile_25__pin_sc_in_0_,
                         left_width_0_height_0_subtile_26__pin_sc_in_0_,
                         left_width_0_height_0_subtile_27__pin_sc_in_0_,
                         left_width_0_height_0_subtile_28__pin_sc_in_0_,
                         left_width_0_height_0_subtile_29__pin_sc_in_0_,
                         left_width_0_height_0_subtile_30__pin_sc_in_0_,
                         left_width_0_height_0_subtile_31__pin_sc_in_0_,
                         left_width_0_height_0_subtile_32__pin_sc_in_0_,
                         left_width_0_height_0_subtile_33__pin_sc_in_0_,
                         left_width_0_height_0_subtile_34__pin_sc_in_0_,
                         left_width_0_height_0_subtile_35__pin_sc_in_0_,
                         left_width_0_height_0_subtile_36__pin_sc_in_0_,
                         left_width_0_height_0_subtile_37__pin_sc_in_0_,
                         left_width_0_height_0_subtile_38__pin_sc_in_0_,
                         left_width_0_height_0_subtile_39__pin_sc_in_0_,
                         left_width_0_height_0_subtile_40__pin_sc_in_0_,
                         left_width_0_height_0_subtile_41__pin_sc_in_0_,
                         left_width_0_height_0_subtile_42__pin_sc_in_0_,
                         left_width_0_height_0_subtile_43__pin_sc_in_0_,
                         left_width_0_height_0_subtile_44__pin_sc_in_0_,
                         left_width_0_height_0_subtile_45__pin_sc_in_0_,
                         left_width_0_height_0_subtile_46__pin_sc_in_0_,
                         left_width_0_height_0_subtile_47__pin_sc_in_0_,
                         left_width_0_height_0_subtile_48__pin_sc_in_0_,
                         left_width_0_height_0_subtile_49__pin_sc_in_0_,
                         left_width_0_height_0_subtile_50__pin_sc_in_0_,
                         left_width_0_height_0_subtile_51__pin_sc_in_0_,
                         left_width_0_height_0_subtile_52__pin_sc_in_0_,
                         left_width_0_height_0_subtile_53__pin_sc_in_0_,
                         left_width_0_height_0_subtile_54__pin_sc_in_0_,
                         left_width_0_height_0_subtile_55__pin_sc_in_0_,
                         left_width_0_height_0_subtile_56__pin_sc_in_0_,
                         left_width_0_height_0_subtile_57__pin_sc_in_0_,
                         left_width_0_height_0_subtile_58__pin_sc_in_0_,
                         left_width_0_height_0_subtile_59__pin_sc_in_0_,
                         ccff_head,
                         top_width_0_height_0_subtile_30__pin_a2f_o_0_,
                         top_width_0_height_0_subtile_30__pin_a2f_o_1_,
                         top_width_0_height_0_subtile_31__pin_a2f_o_0_,
                         top_width_0_height_0_subtile_31__pin_a2f_o_1_,
                         top_width_0_height_0_subtile_32__pin_a2f_o_0_,
                         top_width_0_height_0_subtile_32__pin_a2f_o_1_,
                         top_width_0_height_0_subtile_33__pin_a2f_o_0_,
                         top_width_0_height_0_subtile_33__pin_a2f_o_1_,
                         top_width_0_height_0_subtile_34__pin_a2f_o_0_,
                         top_width_0_height_0_subtile_34__pin_a2f_o_1_,
                         top_width_0_height_0_subtile_35__pin_a2f_o_0_,
                         top_width_0_height_0_subtile_35__pin_a2f_o_1_,
                         top_width_0_height_0_subtile_36__pin_a2f_o_0_,
                         top_width_0_height_0_subtile_36__pin_a2f_o_1_,
                         top_width_0_height_0_subtile_37__pin_a2f_o_0_,
                         top_width_0_height_0_subtile_37__pin_a2f_o_1_,
                         top_width_0_height_0_subtile_38__pin_a2f_o_0_,
                         top_width_0_height_0_subtile_38__pin_a2f_o_1_,
                         top_width_0_height_0_subtile_39__pin_a2f_o_0_,
                         top_width_0_height_0_subtile_39__pin_a2f_o_1_,
                         top_width_0_height_0_subtile_40__pin_a2f_o_0_,
                         top_width_0_height_0_subtile_40__pin_a2f_o_1_,
                         top_width_0_height_0_subtile_41__pin_a2f_o_0_,
                         top_width_0_height_0_subtile_41__pin_a2f_o_1_,
                         top_width_0_height_0_subtile_42__pin_a2f_o_0_,
                         top_width_0_height_0_subtile_42__pin_a2f_o_1_,
                         top_width_0_height_0_subtile_43__pin_a2f_o_0_,
                         top_width_0_height_0_subtile_43__pin_a2f_o_1_,
                         top_width_0_height_0_subtile_44__pin_a2f_o_0_,
                         top_width_0_height_0_subtile_44__pin_a2f_o_1_,
                         top_width_0_height_0_subtile_45__pin_a2f_o_0_,
                         top_width_0_height_0_subtile_45__pin_a2f_o_1_,
                         top_width_0_height_0_subtile_46__pin_a2f_o_0_,
                         top_width_0_height_0_subtile_46__pin_a2f_o_1_,
                         top_width_0_height_0_subtile_47__pin_a2f_o_0_,
                         top_width_0_height_0_subtile_47__pin_a2f_o_1_,
                         top_width_0_height_0_subtile_48__pin_a2f_o_0_,
                         top_width_0_height_0_subtile_48__pin_a2f_o_1_,
                         top_width_0_height_0_subtile_49__pin_a2f_o_0_,
                         top_width_0_height_0_subtile_49__pin_a2f_o_1_,
                         top_width_0_height_0_subtile_50__pin_a2f_o_0_,
                         top_width_0_height_0_subtile_50__pin_a2f_o_1_,
                         top_width_0_height_0_subtile_51__pin_a2f_o_0_,
                         top_width_0_height_0_subtile_51__pin_a2f_o_1_,
                         top_width_0_height_0_subtile_52__pin_a2f_o_0_,
                         top_width_0_height_0_subtile_52__pin_a2f_o_1_,
                         top_width_0_height_0_subtile_53__pin_a2f_o_0_,
                         top_width_0_height_0_subtile_53__pin_a2f_o_1_,
                         top_width_0_height_0_subtile_54__pin_a2f_o_0_,
                         top_width_0_height_0_subtile_54__pin_a2f_o_1_,
                         top_width_0_height_0_subtile_55__pin_a2f_o_0_,
                         top_width_0_height_0_subtile_55__pin_a2f_o_1_,
                         top_width_0_height_0_subtile_56__pin_a2f_o_0_,
                         top_width_0_height_0_subtile_56__pin_a2f_o_1_,
                         top_width_0_height_0_subtile_57__pin_a2f_o_0_,
                         top_width_0_height_0_subtile_57__pin_a2f_o_1_,
                         top_width_0_height_0_subtile_58__pin_a2f_o_0_,
                         top_width_0_height_0_subtile_58__pin_a2f_o_1_,
                         top_width_0_height_0_subtile_59__pin_a2f_o_0_,
                         top_width_0_height_0_subtile_59__pin_a2f_o_1_,
                         right_width_0_height_0_subtile_0__pin_a2f_o_0_,
                         right_width_0_height_0_subtile_0__pin_a2f_o_1_,
                         right_width_0_height_0_subtile_1__pin_a2f_o_0_,
                         right_width_0_height_0_subtile_1__pin_a2f_o_1_,
                         right_width_0_height_0_subtile_2__pin_a2f_o_0_,
                         right_width_0_height_0_subtile_2__pin_a2f_o_1_,
                         right_width_0_height_0_subtile_3__pin_a2f_o_0_,
                         right_width_0_height_0_subtile_3__pin_a2f_o_1_,
                         right_width_0_height_0_subtile_4__pin_a2f_o_0_,
                         right_width_0_height_0_subtile_4__pin_a2f_o_1_,
                         right_width_0_height_0_subtile_5__pin_a2f_o_0_,
                         right_width_0_height_0_subtile_5__pin_a2f_o_1_,
                         right_width_0_height_0_subtile_6__pin_a2f_o_0_,
                         right_width_0_height_0_subtile_6__pin_a2f_o_1_,
                         right_width_0_height_0_subtile_7__pin_a2f_o_0_,
                         right_width_0_height_0_subtile_7__pin_a2f_o_1_,
                         right_width_0_height_0_subtile_8__pin_a2f_o_0_,
                         right_width_0_height_0_subtile_8__pin_a2f_o_1_,
                         right_width_0_height_0_subtile_9__pin_a2f_o_0_,
                         right_width_0_height_0_subtile_9__pin_a2f_o_1_,
                         right_width_0_height_0_subtile_10__pin_a2f_o_0_,
                         right_width_0_height_0_subtile_10__pin_a2f_o_1_,
                         right_width_0_height_0_subtile_11__pin_a2f_o_0_,
                         right_width_0_height_0_subtile_11__pin_a2f_o_1_,
                         right_width_0_height_0_subtile_12__pin_a2f_o_0_,
                         right_width_0_height_0_subtile_12__pin_a2f_o_1_,
                         right_width_0_height_0_subtile_13__pin_a2f_o_0_,
                         right_width_0_height_0_subtile_13__pin_a2f_o_1_,
                         right_width_0_height_0_subtile_14__pin_a2f_o_0_,
                         right_width_0_height_0_subtile_14__pin_a2f_o_1_,
                         right_width_0_height_0_subtile_15__pin_a2f_o_0_,
                         right_width_0_height_0_subtile_15__pin_a2f_o_1_,
                         right_width_0_height_0_subtile_16__pin_a2f_o_0_,
                         right_width_0_height_0_subtile_16__pin_a2f_o_1_,
                         right_width_0_height_0_subtile_17__pin_a2f_o_0_,
                         right_width_0_height_0_subtile_17__pin_a2f_o_1_,
                         right_width_0_height_0_subtile_18__pin_a2f_o_0_,
                         right_width_0_height_0_subtile_18__pin_a2f_o_1_,
                         right_width_0_height_0_subtile_19__pin_a2f_o_0_,
                         right_width_0_height_0_subtile_19__pin_a2f_o_1_,
                         right_width_0_height_0_subtile_20__pin_a2f_o_0_,
                         right_width_0_height_0_subtile_20__pin_a2f_o_1_,
                         right_width_0_height_0_subtile_21__pin_a2f_o_0_,
                         right_width_0_height_0_subtile_21__pin_a2f_o_1_,
                         right_width_0_height_0_subtile_22__pin_a2f_o_0_,
                         right_width_0_height_0_subtile_22__pin_a2f_o_1_,
                         right_width_0_height_0_subtile_23__pin_a2f_o_0_,
                         right_width_0_height_0_subtile_23__pin_a2f_o_1_,
                         right_width_0_height_0_subtile_24__pin_a2f_o_0_,
                         right_width_0_height_0_subtile_24__pin_a2f_o_1_,
                         right_width_0_height_0_subtile_25__pin_a2f_o_0_,
                         right_width_0_height_0_subtile_25__pin_a2f_o_1_,
                         right_width_0_height_0_subtile_26__pin_a2f_o_0_,
                         right_width_0_height_0_subtile_26__pin_a2f_o_1_,
                         right_width_0_height_0_subtile_27__pin_a2f_o_0_,
                         right_width_0_height_0_subtile_27__pin_a2f_o_1_,
                         right_width_0_height_0_subtile_28__pin_a2f_o_0_,
                         right_width_0_height_0_subtile_28__pin_a2f_o_1_,
                         right_width_0_height_0_subtile_29__pin_a2f_o_0_,
                         right_width_0_height_0_subtile_29__pin_a2f_o_1_,
                         left_width_0_height_0_subtile_0__pin_sc_out_0_,
                         left_width_0_height_0_subtile_1__pin_sc_out_0_,
                         left_width_0_height_0_subtile_2__pin_sc_out_0_,
                         left_width_0_height_0_subtile_3__pin_sc_out_0_,
                         left_width_0_height_0_subtile_4__pin_sc_out_0_,
                         left_width_0_height_0_subtile_5__pin_sc_out_0_,
                         left_width_0_height_0_subtile_6__pin_sc_out_0_,
                         left_width_0_height_0_subtile_7__pin_sc_out_0_,
                         left_width_0_height_0_subtile_8__pin_sc_out_0_,
                         left_width_0_height_0_subtile_9__pin_sc_out_0_,
                         left_width_0_height_0_subtile_10__pin_sc_out_0_,
                         left_width_0_height_0_subtile_11__pin_sc_out_0_,
                         left_width_0_height_0_subtile_12__pin_sc_out_0_,
                         left_width_0_height_0_subtile_13__pin_sc_out_0_,
                         left_width_0_height_0_subtile_14__pin_sc_out_0_,
                         left_width_0_height_0_subtile_15__pin_sc_out_0_,
                         left_width_0_height_0_subtile_16__pin_sc_out_0_,
                         left_width_0_height_0_subtile_17__pin_sc_out_0_,
                         left_width_0_height_0_subtile_18__pin_sc_out_0_,
                         left_width_0_height_0_subtile_19__pin_sc_out_0_,
                         left_width_0_height_0_subtile_20__pin_sc_out_0_,
                         left_width_0_height_0_subtile_21__pin_sc_out_0_,
                         left_width_0_height_0_subtile_22__pin_sc_out_0_,
                         left_width_0_height_0_subtile_23__pin_sc_out_0_,
                         left_width_0_height_0_subtile_24__pin_sc_out_0_,
                         left_width_0_height_0_subtile_25__pin_sc_out_0_,
                         left_width_0_height_0_subtile_26__pin_sc_out_0_,
                         left_width_0_height_0_subtile_27__pin_sc_out_0_,
                         left_width_0_height_0_subtile_28__pin_sc_out_0_,
                         left_width_0_height_0_subtile_29__pin_sc_out_0_,
                         left_width_0_height_0_subtile_30__pin_sc_out_0_,
                         left_width_0_height_0_subtile_31__pin_sc_out_0_,
                         left_width_0_height_0_subtile_32__pin_sc_out_0_,
                         left_width_0_height_0_subtile_33__pin_sc_out_0_,
                         left_width_0_height_0_subtile_34__pin_sc_out_0_,
                         left_width_0_height_0_subtile_35__pin_sc_out_0_,
                         left_width_0_height_0_subtile_36__pin_sc_out_0_,
                         left_width_0_height_0_subtile_37__pin_sc_out_0_,
                         left_width_0_height_0_subtile_38__pin_sc_out_0_,
                         left_width_0_height_0_subtile_39__pin_sc_out_0_,
                         left_width_0_height_0_subtile_40__pin_sc_out_0_,
                         left_width_0_height_0_subtile_41__pin_sc_out_0_,
                         left_width_0_height_0_subtile_42__pin_sc_out_0_,
                         left_width_0_height_0_subtile_43__pin_sc_out_0_,
                         left_width_0_height_0_subtile_44__pin_sc_out_0_,
                         left_width_0_height_0_subtile_45__pin_sc_out_0_,
                         left_width_0_height_0_subtile_46__pin_sc_out_0_,
                         left_width_0_height_0_subtile_47__pin_sc_out_0_,
                         left_width_0_height_0_subtile_48__pin_sc_out_0_,
                         left_width_0_height_0_subtile_49__pin_sc_out_0_,
                         left_width_0_height_0_subtile_50__pin_sc_out_0_,
                         left_width_0_height_0_subtile_51__pin_sc_out_0_,
                         left_width_0_height_0_subtile_52__pin_sc_out_0_,
                         left_width_0_height_0_subtile_53__pin_sc_out_0_,
                         left_width_0_height_0_subtile_54__pin_sc_out_0_,
                         left_width_0_height_0_subtile_55__pin_sc_out_0_,
                         left_width_0_height_0_subtile_56__pin_sc_out_0_,
                         left_width_0_height_0_subtile_57__pin_sc_out_0_,
                         left_width_0_height_0_subtile_58__pin_sc_out_0_,
                         left_width_0_height_0_subtile_59__pin_sc_out_0_,
                         ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] global_reset;
//----- GLOBAL PORTS -----
input [0:0] scan_mode;
//----- GLOBAL PORTS -----
input [0:0] scan_enable;
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_clock;
//----- GPIN PORTS -----
input [0:59] gfpga_pad_RS_PREIO_A2F;
//----- GPOUT PORTS -----
output [0:59] gfpga_pad_RS_PREIO_F2A;
//----- GPOUT PORTS -----
output [0:59] gfpga_pad_RS_PREIO_SOC_CLK;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_14__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_15__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_16__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_17__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_18__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_19__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_20__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_21__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_22__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_23__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_24__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_25__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_26__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_27__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_28__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_29__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_30__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_31__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_32__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_33__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_34__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_35__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_36__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_37__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_38__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_39__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_40__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_41__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_42__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_43__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_44__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_45__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_46__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_47__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_48__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_49__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_50__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_51__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_52__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_53__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_54__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_55__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_56__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_57__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_58__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_59__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_1__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_2__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_3__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_4__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_5__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_6__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_7__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_8__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_9__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_10__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_11__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_12__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_13__pin_f2a_i_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_1__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_1__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_1__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_1__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_1__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_1__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_1__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_1__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_1__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_1__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_1__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_1__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_1__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_1__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_1__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_1__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_2__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_2__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_2__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_2__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_2__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_2__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_2__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_2__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_2__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_2__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_2__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_2__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_2__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_2__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_2__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_2__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_3__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_3__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_3__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_3__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_3__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_3__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_3__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_3__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_3__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_3__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_3__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_3__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_3__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_3__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_3__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_3__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_4__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_4__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_4__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_4__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_4__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_4__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_4__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_4__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_4__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_4__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_4__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_4__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_4__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_4__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_4__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_4__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_5__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_5__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_5__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_5__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_5__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_5__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_5__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_5__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_5__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_5__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_5__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_5__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_5__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_5__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_5__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_5__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_6__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_6__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_6__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_6__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_6__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_6__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_6__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_6__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_6__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_6__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_6__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_6__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_6__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_6__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_6__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_6__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_7__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_7__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_7__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_7__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_7__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_7__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_7__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_7__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_7__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_7__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_7__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_7__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_7__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_7__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_7__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_7__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_8__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_8__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_8__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_8__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_8__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_8__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_8__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_8__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_8__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_8__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_8__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_8__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_8__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_8__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_8__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_8__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_9__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_9__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_9__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_9__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_9__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_9__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_9__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_9__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_9__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_9__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_9__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_9__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_9__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_9__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_9__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_9__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_10__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_10__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_10__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_10__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_10__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_10__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_10__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_10__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_10__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_10__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_10__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_10__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_10__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_10__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_10__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_10__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_11__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_11__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_11__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_11__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_11__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_11__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_11__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_11__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_11__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_11__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_11__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_11__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_11__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_11__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_11__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_11__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_12__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_12__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_12__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_12__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_12__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_12__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_12__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_12__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_12__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_12__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_12__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_12__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_12__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_12__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_12__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_12__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_13__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_13__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_13__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_13__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_13__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_13__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_13__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_13__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_13__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_13__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_13__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_13__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_13__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_13__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_13__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_13__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_14__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_14__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_14__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_14__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_14__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_14__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_14__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_14__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_14__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_14__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_14__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_14__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_14__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_14__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_14__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_14__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_15__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_15__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_15__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_15__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_15__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_15__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_15__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_15__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_15__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_15__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_15__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_15__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_15__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_15__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_15__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_15__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_16__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_16__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_16__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_16__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_16__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_16__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_16__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_16__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_16__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_16__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_16__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_16__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_16__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_16__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_16__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_16__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_17__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_17__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_17__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_17__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_17__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_17__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_17__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_17__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_17__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_17__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_17__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_17__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_17__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_17__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_17__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_17__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_18__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_18__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_18__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_18__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_18__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_18__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_18__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_18__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_18__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_18__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_18__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_18__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_18__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_18__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_18__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_18__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_19__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_19__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_19__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_19__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_19__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_19__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_19__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_19__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_19__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_19__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_19__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_19__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_19__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_19__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_19__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_19__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_20__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_20__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_20__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_20__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_20__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_20__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_20__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_20__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_20__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_20__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_20__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_20__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_20__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_20__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_20__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_20__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_21__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_21__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_21__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_21__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_21__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_21__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_21__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_21__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_21__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_21__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_21__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_21__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_21__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_21__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_21__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_21__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_22__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_22__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_22__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_22__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_22__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_22__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_22__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_22__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_22__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_22__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_22__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_22__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_22__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_22__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_22__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_22__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_23__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_23__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_23__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_23__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_23__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_23__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_23__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_23__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_23__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_23__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_23__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_23__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_23__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_23__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_23__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_23__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_24__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_24__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_24__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_24__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_24__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_24__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_24__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_24__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_24__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_24__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_24__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_24__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_24__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_24__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_24__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_24__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_25__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_25__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_25__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_25__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_25__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_25__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_25__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_25__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_25__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_25__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_25__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_25__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_25__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_25__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_25__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_25__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_26__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_26__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_26__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_26__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_26__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_26__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_26__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_26__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_26__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_26__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_26__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_26__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_26__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_26__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_26__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_26__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_27__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_27__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_27__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_27__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_27__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_27__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_27__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_27__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_27__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_27__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_27__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_27__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_27__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_27__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_27__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_27__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_28__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_28__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_28__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_28__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_28__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_28__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_28__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_28__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_28__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_28__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_28__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_28__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_28__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_28__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_28__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_28__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_29__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_29__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_29__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_29__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_29__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_29__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_29__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_29__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_29__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_29__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_29__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_29__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_29__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_29__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_29__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_29__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_30__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_30__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_30__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_30__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_30__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_30__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_30__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_30__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_30__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_30__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_30__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_30__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_30__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_30__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_30__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_30__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_31__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_31__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_31__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_31__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_31__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_31__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_31__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_31__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_31__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_31__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_31__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_31__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_31__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_31__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_31__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_31__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_32__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_32__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_32__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_32__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_32__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_32__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_32__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_32__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_32__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_32__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_32__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_32__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_32__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_32__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_32__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_32__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_33__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_33__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_33__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_33__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_33__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_33__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_33__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_33__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_33__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_33__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_33__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_33__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_33__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_33__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_33__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_33__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_34__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_34__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_34__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_34__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_34__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_34__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_34__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_34__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_34__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_34__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_34__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_34__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_34__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_34__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_34__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_34__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_35__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_35__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_35__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_35__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_35__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_35__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_35__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_35__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_35__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_35__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_35__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_35__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_35__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_35__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_35__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_35__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_36__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_36__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_36__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_36__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_36__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_36__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_36__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_36__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_36__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_36__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_36__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_36__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_36__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_36__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_36__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_36__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_37__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_37__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_37__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_37__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_37__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_37__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_37__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_37__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_37__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_37__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_37__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_37__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_37__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_37__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_37__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_37__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_38__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_38__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_38__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_38__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_38__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_38__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_38__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_38__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_38__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_38__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_38__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_38__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_38__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_38__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_38__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_38__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_39__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_39__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_39__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_39__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_39__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_39__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_39__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_39__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_39__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_39__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_39__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_39__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_39__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_39__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_39__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_39__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_40__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_40__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_40__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_40__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_40__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_40__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_40__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_40__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_40__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_40__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_40__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_40__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_40__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_40__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_40__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_40__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_41__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_41__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_41__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_41__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_41__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_41__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_41__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_41__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_41__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_41__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_41__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_41__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_41__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_41__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_41__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_41__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_42__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_42__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_42__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_42__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_42__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_42__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_42__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_42__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_42__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_42__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_42__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_42__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_42__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_42__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_42__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_42__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_43__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_43__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_43__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_43__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_43__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_43__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_43__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_43__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_43__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_43__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_43__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_43__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_43__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_43__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_43__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_43__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_44__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_44__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_44__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_44__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_44__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_44__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_44__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_44__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_44__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_44__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_44__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_44__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_44__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_44__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_44__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_44__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_45__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_45__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_45__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_45__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_45__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_45__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_45__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_45__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_45__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_45__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_45__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_45__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_45__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_45__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_45__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_45__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_46__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_46__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_46__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_46__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_46__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_46__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_46__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_46__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_46__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_46__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_46__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_46__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_46__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_46__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_46__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_46__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_47__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_47__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_47__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_47__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_47__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_47__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_47__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_47__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_47__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_47__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_47__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_47__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_47__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_47__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_47__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_47__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_48__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_48__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_48__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_48__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_48__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_48__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_48__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_48__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_48__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_48__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_48__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_48__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_48__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_48__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_48__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_48__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_49__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_49__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_49__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_49__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_49__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_49__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_49__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_49__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_49__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_49__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_49__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_49__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_49__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_49__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_49__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_49__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_50__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_50__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_50__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_50__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_50__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_50__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_50__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_50__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_50__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_50__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_50__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_50__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_50__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_50__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_50__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_50__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_51__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_51__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_51__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_51__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_51__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_51__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_51__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_51__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_51__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_51__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_51__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_51__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_51__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_51__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_51__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_51__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_52__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_52__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_52__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_52__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_52__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_52__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_52__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_52__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_52__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_52__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_52__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_52__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_52__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_52__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_52__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_52__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_53__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_53__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_53__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_53__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_53__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_53__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_53__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_53__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_53__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_53__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_53__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_53__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_53__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_53__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_53__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_53__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_54__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_54__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_54__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_54__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_54__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_54__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_54__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_54__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_54__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_54__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_54__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_54__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_54__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_54__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_54__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_54__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_55__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_55__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_55__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_55__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_55__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_55__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_55__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_55__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_55__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_55__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_55__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_55__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_55__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_55__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_55__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_55__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_56__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_56__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_56__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_56__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_56__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_56__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_56__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_56__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_56__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_56__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_56__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_56__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_56__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_56__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_56__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_56__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_57__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_57__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_57__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_57__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_57__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_57__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_57__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_57__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_57__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_57__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_57__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_57__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_57__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_57__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_57__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_57__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_58__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_58__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_58__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_58__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_58__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_58__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_58__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_58__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_58__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_58__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_58__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_58__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_58__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_58__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_58__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_58__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_59__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_59__pin_clk_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_59__pin_clk_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_59__pin_clk_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_59__pin_clk_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_59__pin_clk_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_59__pin_clk_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_59__pin_clk_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_59__pin_clk_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_59__pin_clk_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_59__pin_clk_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_59__pin_clk_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_59__pin_clk_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_59__pin_clk_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_59__pin_clk_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_59__pin_clk_15_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_1__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_2__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_3__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_4__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_5__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_6__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_7__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_8__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_9__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_10__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_11__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_12__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_13__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_14__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_15__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_16__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_17__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_18__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_19__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_20__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_21__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_22__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_23__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_24__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_25__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_26__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_27__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_28__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_29__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_30__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_31__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_32__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_33__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_34__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_35__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_36__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_37__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_38__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_39__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_40__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_41__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_42__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_43__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_44__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_45__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_46__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_47__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_48__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_49__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_50__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_51__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_52__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_53__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_54__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_55__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_56__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_57__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_58__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_59__pin_sc_in_0_;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_30__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_30__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_31__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_31__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_32__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_32__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_33__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_33__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_34__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_34__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_35__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_35__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_36__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_36__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_37__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_37__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_38__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_38__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_39__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_39__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_40__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_40__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_41__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_41__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_42__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_42__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_43__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_43__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_44__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_44__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_45__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_45__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_46__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_46__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_47__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_47__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_48__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_48__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_49__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_49__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_50__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_50__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_51__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_51__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_52__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_52__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_53__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_53__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_54__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_54__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_55__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_55__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_56__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_56__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_57__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_57__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_58__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_58__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_59__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_59__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_1__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_1__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_2__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_2__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_3__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_3__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_4__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_4__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_5__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_5__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_6__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_6__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_7__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_7__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_8__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_8__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_9__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_9__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_10__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_10__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_11__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_11__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_12__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_12__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_13__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_13__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_14__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_14__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_15__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_15__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_16__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_16__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_17__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_17__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_18__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_18__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_19__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_19__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_20__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_20__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_21__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_21__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_22__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_22__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_23__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_23__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_24__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_24__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_25__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_25__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_26__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_26__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_27__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_27__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_28__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_28__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_29__pin_a2f_o_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_29__pin_a2f_o_1_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_1__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_2__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_3__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_4__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_5__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_6__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_7__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_8__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_9__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_10__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_11__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_12__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_13__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_14__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_15__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_16__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_17__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_18__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_19__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_20__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_21__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_22__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_23__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_24__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_25__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_26__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_27__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_28__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_29__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_30__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_31__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_32__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_33__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_34__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_35__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_36__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_37__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_38__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_39__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_40__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_41__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_42__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_43__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_44__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_45__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_46__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_47__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_48__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_49__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_50__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_51__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_52__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_53__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_54__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_55__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_56__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_57__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_58__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_59__pin_sc_out_0_;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__0 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[0]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[0]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[0]),
		.io_corner_f2a_i(right_width_0_height_0_subtile_0__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_0__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_0__pin_clk_0_, bottom_width_0_height_0_subtile_0__pin_clk_1_, bottom_width_0_height_0_subtile_0__pin_clk_2_, bottom_width_0_height_0_subtile_0__pin_clk_3_, bottom_width_0_height_0_subtile_0__pin_clk_4_, bottom_width_0_height_0_subtile_0__pin_clk_5_, bottom_width_0_height_0_subtile_0__pin_clk_6_, bottom_width_0_height_0_subtile_0__pin_clk_7_, bottom_width_0_height_0_subtile_0__pin_clk_8_, bottom_width_0_height_0_subtile_0__pin_clk_9_, bottom_width_0_height_0_subtile_0__pin_clk_10_, bottom_width_0_height_0_subtile_0__pin_clk_11_, bottom_width_0_height_0_subtile_0__pin_clk_12_, bottom_width_0_height_0_subtile_0__pin_clk_13_, bottom_width_0_height_0_subtile_0__pin_clk_14_, bottom_width_0_height_0_subtile_0__pin_clk_15_}),
		.ccff_head(ccff_head),
		.io_corner_a2f_o({right_width_0_height_0_subtile_0__pin_a2f_o_0_, right_width_0_height_0_subtile_0__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_0__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_corner_mode_io_corner__0_ccff_tail));

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__1 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[1]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[1]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[1]),
		.io_corner_f2a_i(right_width_0_height_0_subtile_1__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_1__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_1__pin_clk_0_, bottom_width_0_height_0_subtile_1__pin_clk_1_, bottom_width_0_height_0_subtile_1__pin_clk_2_, bottom_width_0_height_0_subtile_1__pin_clk_3_, bottom_width_0_height_0_subtile_1__pin_clk_4_, bottom_width_0_height_0_subtile_1__pin_clk_5_, bottom_width_0_height_0_subtile_1__pin_clk_6_, bottom_width_0_height_0_subtile_1__pin_clk_7_, bottom_width_0_height_0_subtile_1__pin_clk_8_, bottom_width_0_height_0_subtile_1__pin_clk_9_, bottom_width_0_height_0_subtile_1__pin_clk_10_, bottom_width_0_height_0_subtile_1__pin_clk_11_, bottom_width_0_height_0_subtile_1__pin_clk_12_, bottom_width_0_height_0_subtile_1__pin_clk_13_, bottom_width_0_height_0_subtile_1__pin_clk_14_, bottom_width_0_height_0_subtile_1__pin_clk_15_}),
		.ccff_head(logical_tile_io_corner_mode_io_corner__0_ccff_tail),
		.io_corner_a2f_o({right_width_0_height_0_subtile_1__pin_a2f_o_0_, right_width_0_height_0_subtile_1__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_1__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_corner_mode_io_corner__1_ccff_tail));

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__2 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[2]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[2]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[2]),
		.io_corner_f2a_i(right_width_0_height_0_subtile_2__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_2__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_2__pin_clk_0_, bottom_width_0_height_0_subtile_2__pin_clk_1_, bottom_width_0_height_0_subtile_2__pin_clk_2_, bottom_width_0_height_0_subtile_2__pin_clk_3_, bottom_width_0_height_0_subtile_2__pin_clk_4_, bottom_width_0_height_0_subtile_2__pin_clk_5_, bottom_width_0_height_0_subtile_2__pin_clk_6_, bottom_width_0_height_0_subtile_2__pin_clk_7_, bottom_width_0_height_0_subtile_2__pin_clk_8_, bottom_width_0_height_0_subtile_2__pin_clk_9_, bottom_width_0_height_0_subtile_2__pin_clk_10_, bottom_width_0_height_0_subtile_2__pin_clk_11_, bottom_width_0_height_0_subtile_2__pin_clk_12_, bottom_width_0_height_0_subtile_2__pin_clk_13_, bottom_width_0_height_0_subtile_2__pin_clk_14_, bottom_width_0_height_0_subtile_2__pin_clk_15_}),
		.ccff_head(logical_tile_io_corner_mode_io_corner__1_ccff_tail),
		.io_corner_a2f_o({right_width_0_height_0_subtile_2__pin_a2f_o_0_, right_width_0_height_0_subtile_2__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_2__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_corner_mode_io_corner__2_ccff_tail));

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__3 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[3]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[3]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[3]),
		.io_corner_f2a_i(right_width_0_height_0_subtile_3__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_3__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_3__pin_clk_0_, bottom_width_0_height_0_subtile_3__pin_clk_1_, bottom_width_0_height_0_subtile_3__pin_clk_2_, bottom_width_0_height_0_subtile_3__pin_clk_3_, bottom_width_0_height_0_subtile_3__pin_clk_4_, bottom_width_0_height_0_subtile_3__pin_clk_5_, bottom_width_0_height_0_subtile_3__pin_clk_6_, bottom_width_0_height_0_subtile_3__pin_clk_7_, bottom_width_0_height_0_subtile_3__pin_clk_8_, bottom_width_0_height_0_subtile_3__pin_clk_9_, bottom_width_0_height_0_subtile_3__pin_clk_10_, bottom_width_0_height_0_subtile_3__pin_clk_11_, bottom_width_0_height_0_subtile_3__pin_clk_12_, bottom_width_0_height_0_subtile_3__pin_clk_13_, bottom_width_0_height_0_subtile_3__pin_clk_14_, bottom_width_0_height_0_subtile_3__pin_clk_15_}),
		.ccff_head(logical_tile_io_corner_mode_io_corner__2_ccff_tail),
		.io_corner_a2f_o({right_width_0_height_0_subtile_3__pin_a2f_o_0_, right_width_0_height_0_subtile_3__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_3__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_corner_mode_io_corner__3_ccff_tail));

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__4 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[4]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[4]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[4]),
		.io_corner_f2a_i(right_width_0_height_0_subtile_4__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_4__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_4__pin_clk_0_, bottom_width_0_height_0_subtile_4__pin_clk_1_, bottom_width_0_height_0_subtile_4__pin_clk_2_, bottom_width_0_height_0_subtile_4__pin_clk_3_, bottom_width_0_height_0_subtile_4__pin_clk_4_, bottom_width_0_height_0_subtile_4__pin_clk_5_, bottom_width_0_height_0_subtile_4__pin_clk_6_, bottom_width_0_height_0_subtile_4__pin_clk_7_, bottom_width_0_height_0_subtile_4__pin_clk_8_, bottom_width_0_height_0_subtile_4__pin_clk_9_, bottom_width_0_height_0_subtile_4__pin_clk_10_, bottom_width_0_height_0_subtile_4__pin_clk_11_, bottom_width_0_height_0_subtile_4__pin_clk_12_, bottom_width_0_height_0_subtile_4__pin_clk_13_, bottom_width_0_height_0_subtile_4__pin_clk_14_, bottom_width_0_height_0_subtile_4__pin_clk_15_}),
		.ccff_head(logical_tile_io_corner_mode_io_corner__3_ccff_tail),
		.io_corner_a2f_o({right_width_0_height_0_subtile_4__pin_a2f_o_0_, right_width_0_height_0_subtile_4__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_4__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_corner_mode_io_corner__4_ccff_tail));

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__5 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[5]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[5]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[5]),
		.io_corner_f2a_i(right_width_0_height_0_subtile_5__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_5__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_5__pin_clk_0_, bottom_width_0_height_0_subtile_5__pin_clk_1_, bottom_width_0_height_0_subtile_5__pin_clk_2_, bottom_width_0_height_0_subtile_5__pin_clk_3_, bottom_width_0_height_0_subtile_5__pin_clk_4_, bottom_width_0_height_0_subtile_5__pin_clk_5_, bottom_width_0_height_0_subtile_5__pin_clk_6_, bottom_width_0_height_0_subtile_5__pin_clk_7_, bottom_width_0_height_0_subtile_5__pin_clk_8_, bottom_width_0_height_0_subtile_5__pin_clk_9_, bottom_width_0_height_0_subtile_5__pin_clk_10_, bottom_width_0_height_0_subtile_5__pin_clk_11_, bottom_width_0_height_0_subtile_5__pin_clk_12_, bottom_width_0_height_0_subtile_5__pin_clk_13_, bottom_width_0_height_0_subtile_5__pin_clk_14_, bottom_width_0_height_0_subtile_5__pin_clk_15_}),
		.ccff_head(logical_tile_io_corner_mode_io_corner__4_ccff_tail),
		.io_corner_a2f_o({right_width_0_height_0_subtile_5__pin_a2f_o_0_, right_width_0_height_0_subtile_5__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_5__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_corner_mode_io_corner__5_ccff_tail));

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__6 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[6]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[6]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[6]),
		.io_corner_f2a_i(right_width_0_height_0_subtile_6__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_6__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_6__pin_clk_0_, bottom_width_0_height_0_subtile_6__pin_clk_1_, bottom_width_0_height_0_subtile_6__pin_clk_2_, bottom_width_0_height_0_subtile_6__pin_clk_3_, bottom_width_0_height_0_subtile_6__pin_clk_4_, bottom_width_0_height_0_subtile_6__pin_clk_5_, bottom_width_0_height_0_subtile_6__pin_clk_6_, bottom_width_0_height_0_subtile_6__pin_clk_7_, bottom_width_0_height_0_subtile_6__pin_clk_8_, bottom_width_0_height_0_subtile_6__pin_clk_9_, bottom_width_0_height_0_subtile_6__pin_clk_10_, bottom_width_0_height_0_subtile_6__pin_clk_11_, bottom_width_0_height_0_subtile_6__pin_clk_12_, bottom_width_0_height_0_subtile_6__pin_clk_13_, bottom_width_0_height_0_subtile_6__pin_clk_14_, bottom_width_0_height_0_subtile_6__pin_clk_15_}),
		.ccff_head(logical_tile_io_corner_mode_io_corner__5_ccff_tail),
		.io_corner_a2f_o({right_width_0_height_0_subtile_6__pin_a2f_o_0_, right_width_0_height_0_subtile_6__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_6__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_corner_mode_io_corner__6_ccff_tail));

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__7 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[7]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[7]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[7]),
		.io_corner_f2a_i(right_width_0_height_0_subtile_7__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_7__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_7__pin_clk_0_, bottom_width_0_height_0_subtile_7__pin_clk_1_, bottom_width_0_height_0_subtile_7__pin_clk_2_, bottom_width_0_height_0_subtile_7__pin_clk_3_, bottom_width_0_height_0_subtile_7__pin_clk_4_, bottom_width_0_height_0_subtile_7__pin_clk_5_, bottom_width_0_height_0_subtile_7__pin_clk_6_, bottom_width_0_height_0_subtile_7__pin_clk_7_, bottom_width_0_height_0_subtile_7__pin_clk_8_, bottom_width_0_height_0_subtile_7__pin_clk_9_, bottom_width_0_height_0_subtile_7__pin_clk_10_, bottom_width_0_height_0_subtile_7__pin_clk_11_, bottom_width_0_height_0_subtile_7__pin_clk_12_, bottom_width_0_height_0_subtile_7__pin_clk_13_, bottom_width_0_height_0_subtile_7__pin_clk_14_, bottom_width_0_height_0_subtile_7__pin_clk_15_}),
		.ccff_head(logical_tile_io_corner_mode_io_corner__6_ccff_tail),
		.io_corner_a2f_o({right_width_0_height_0_subtile_7__pin_a2f_o_0_, right_width_0_height_0_subtile_7__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_7__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_corner_mode_io_corner__7_ccff_tail));

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__8 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[8]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[8]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[8]),
		.io_corner_f2a_i(right_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_8__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_8__pin_clk_0_, bottom_width_0_height_0_subtile_8__pin_clk_1_, bottom_width_0_height_0_subtile_8__pin_clk_2_, bottom_width_0_height_0_subtile_8__pin_clk_3_, bottom_width_0_height_0_subtile_8__pin_clk_4_, bottom_width_0_height_0_subtile_8__pin_clk_5_, bottom_width_0_height_0_subtile_8__pin_clk_6_, bottom_width_0_height_0_subtile_8__pin_clk_7_, bottom_width_0_height_0_subtile_8__pin_clk_8_, bottom_width_0_height_0_subtile_8__pin_clk_9_, bottom_width_0_height_0_subtile_8__pin_clk_10_, bottom_width_0_height_0_subtile_8__pin_clk_11_, bottom_width_0_height_0_subtile_8__pin_clk_12_, bottom_width_0_height_0_subtile_8__pin_clk_13_, bottom_width_0_height_0_subtile_8__pin_clk_14_, bottom_width_0_height_0_subtile_8__pin_clk_15_}),
		.ccff_head(logical_tile_io_corner_mode_io_corner__7_ccff_tail),
		.io_corner_a2f_o({right_width_0_height_0_subtile_8__pin_a2f_o_0_, right_width_0_height_0_subtile_8__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_8__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_corner_mode_io_corner__8_ccff_tail));

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__9 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[9]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[9]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[9]),
		.io_corner_f2a_i(right_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_9__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_9__pin_clk_0_, bottom_width_0_height_0_subtile_9__pin_clk_1_, bottom_width_0_height_0_subtile_9__pin_clk_2_, bottom_width_0_height_0_subtile_9__pin_clk_3_, bottom_width_0_height_0_subtile_9__pin_clk_4_, bottom_width_0_height_0_subtile_9__pin_clk_5_, bottom_width_0_height_0_subtile_9__pin_clk_6_, bottom_width_0_height_0_subtile_9__pin_clk_7_, bottom_width_0_height_0_subtile_9__pin_clk_8_, bottom_width_0_height_0_subtile_9__pin_clk_9_, bottom_width_0_height_0_subtile_9__pin_clk_10_, bottom_width_0_height_0_subtile_9__pin_clk_11_, bottom_width_0_height_0_subtile_9__pin_clk_12_, bottom_width_0_height_0_subtile_9__pin_clk_13_, bottom_width_0_height_0_subtile_9__pin_clk_14_, bottom_width_0_height_0_subtile_9__pin_clk_15_}),
		.ccff_head(logical_tile_io_corner_mode_io_corner__8_ccff_tail),
		.io_corner_a2f_o({right_width_0_height_0_subtile_9__pin_a2f_o_0_, right_width_0_height_0_subtile_9__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_9__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_corner_mode_io_corner__9_ccff_tail));

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__10 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[10]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[10]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[10]),
		.io_corner_f2a_i(right_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_10__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_10__pin_clk_0_, bottom_width_0_height_0_subtile_10__pin_clk_1_, bottom_width_0_height_0_subtile_10__pin_clk_2_, bottom_width_0_height_0_subtile_10__pin_clk_3_, bottom_width_0_height_0_subtile_10__pin_clk_4_, bottom_width_0_height_0_subtile_10__pin_clk_5_, bottom_width_0_height_0_subtile_10__pin_clk_6_, bottom_width_0_height_0_subtile_10__pin_clk_7_, bottom_width_0_height_0_subtile_10__pin_clk_8_, bottom_width_0_height_0_subtile_10__pin_clk_9_, bottom_width_0_height_0_subtile_10__pin_clk_10_, bottom_width_0_height_0_subtile_10__pin_clk_11_, bottom_width_0_height_0_subtile_10__pin_clk_12_, bottom_width_0_height_0_subtile_10__pin_clk_13_, bottom_width_0_height_0_subtile_10__pin_clk_14_, bottom_width_0_height_0_subtile_10__pin_clk_15_}),
		.ccff_head(logical_tile_io_corner_mode_io_corner__9_ccff_tail),
		.io_corner_a2f_o({right_width_0_height_0_subtile_10__pin_a2f_o_0_, right_width_0_height_0_subtile_10__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_10__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_corner_mode_io_corner__10_ccff_tail));

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__11 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[11]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[11]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[11]),
		.io_corner_f2a_i(right_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_11__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_11__pin_clk_0_, bottom_width_0_height_0_subtile_11__pin_clk_1_, bottom_width_0_height_0_subtile_11__pin_clk_2_, bottom_width_0_height_0_subtile_11__pin_clk_3_, bottom_width_0_height_0_subtile_11__pin_clk_4_, bottom_width_0_height_0_subtile_11__pin_clk_5_, bottom_width_0_height_0_subtile_11__pin_clk_6_, bottom_width_0_height_0_subtile_11__pin_clk_7_, bottom_width_0_height_0_subtile_11__pin_clk_8_, bottom_width_0_height_0_subtile_11__pin_clk_9_, bottom_width_0_height_0_subtile_11__pin_clk_10_, bottom_width_0_height_0_subtile_11__pin_clk_11_, bottom_width_0_height_0_subtile_11__pin_clk_12_, bottom_width_0_height_0_subtile_11__pin_clk_13_, bottom_width_0_height_0_subtile_11__pin_clk_14_, bottom_width_0_height_0_subtile_11__pin_clk_15_}),
		.ccff_head(logical_tile_io_corner_mode_io_corner__10_ccff_tail),
		.io_corner_a2f_o({right_width_0_height_0_subtile_11__pin_a2f_o_0_, right_width_0_height_0_subtile_11__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_11__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_corner_mode_io_corner__11_ccff_tail));

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__12 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[12]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[12]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[12]),
		.io_corner_f2a_i(right_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_12__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_12__pin_clk_0_, bottom_width_0_height_0_subtile_12__pin_clk_1_, bottom_width_0_height_0_subtile_12__pin_clk_2_, bottom_width_0_height_0_subtile_12__pin_clk_3_, bottom_width_0_height_0_subtile_12__pin_clk_4_, bottom_width_0_height_0_subtile_12__pin_clk_5_, bottom_width_0_height_0_subtile_12__pin_clk_6_, bottom_width_0_height_0_subtile_12__pin_clk_7_, bottom_width_0_height_0_subtile_12__pin_clk_8_, bottom_width_0_height_0_subtile_12__pin_clk_9_, bottom_width_0_height_0_subtile_12__pin_clk_10_, bottom_width_0_height_0_subtile_12__pin_clk_11_, bottom_width_0_height_0_subtile_12__pin_clk_12_, bottom_width_0_height_0_subtile_12__pin_clk_13_, bottom_width_0_height_0_subtile_12__pin_clk_14_, bottom_width_0_height_0_subtile_12__pin_clk_15_}),
		.ccff_head(logical_tile_io_corner_mode_io_corner__11_ccff_tail),
		.io_corner_a2f_o({right_width_0_height_0_subtile_12__pin_a2f_o_0_, right_width_0_height_0_subtile_12__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_12__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_corner_mode_io_corner__12_ccff_tail));

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__13 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[13]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[13]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[13]),
		.io_corner_f2a_i(right_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_13__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_13__pin_clk_0_, bottom_width_0_height_0_subtile_13__pin_clk_1_, bottom_width_0_height_0_subtile_13__pin_clk_2_, bottom_width_0_height_0_subtile_13__pin_clk_3_, bottom_width_0_height_0_subtile_13__pin_clk_4_, bottom_width_0_height_0_subtile_13__pin_clk_5_, bottom_width_0_height_0_subtile_13__pin_clk_6_, bottom_width_0_height_0_subtile_13__pin_clk_7_, bottom_width_0_height_0_subtile_13__pin_clk_8_, bottom_width_0_height_0_subtile_13__pin_clk_9_, bottom_width_0_height_0_subtile_13__pin_clk_10_, bottom_width_0_height_0_subtile_13__pin_clk_11_, bottom_width_0_height_0_subtile_13__pin_clk_12_, bottom_width_0_height_0_subtile_13__pin_clk_13_, bottom_width_0_height_0_subtile_13__pin_clk_14_, bottom_width_0_height_0_subtile_13__pin_clk_15_}),
		.ccff_head(logical_tile_io_corner_mode_io_corner__12_ccff_tail),
		.io_corner_a2f_o({right_width_0_height_0_subtile_13__pin_a2f_o_0_, right_width_0_height_0_subtile_13__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_13__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_corner_mode_io_corner__13_ccff_tail));

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__14 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[14]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[14]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[14]),
		.io_corner_f2a_i(top_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_14__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_14__pin_clk_0_, bottom_width_0_height_0_subtile_14__pin_clk_1_, bottom_width_0_height_0_subtile_14__pin_clk_2_, bottom_width_0_height_0_subtile_14__pin_clk_3_, bottom_width_0_height_0_subtile_14__pin_clk_4_, bottom_width_0_height_0_subtile_14__pin_clk_5_, bottom_width_0_height_0_subtile_14__pin_clk_6_, bottom_width_0_height_0_subtile_14__pin_clk_7_, bottom_width_0_height_0_subtile_14__pin_clk_8_, bottom_width_0_height_0_subtile_14__pin_clk_9_, bottom_width_0_height_0_subtile_14__pin_clk_10_, bottom_width_0_height_0_subtile_14__pin_clk_11_, bottom_width_0_height_0_subtile_14__pin_clk_12_, bottom_width_0_height_0_subtile_14__pin_clk_13_, bottom_width_0_height_0_subtile_14__pin_clk_14_, bottom_width_0_height_0_subtile_14__pin_clk_15_}),
		.ccff_head(logical_tile_io_corner_mode_io_corner__13_ccff_tail),
		.io_corner_a2f_o({right_width_0_height_0_subtile_14__pin_a2f_o_0_, right_width_0_height_0_subtile_14__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_14__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_corner_mode_io_corner__14_ccff_tail));

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__15 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[15]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[15]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[15]),
		.io_corner_f2a_i(top_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_15__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_15__pin_clk_0_, bottom_width_0_height_0_subtile_15__pin_clk_1_, bottom_width_0_height_0_subtile_15__pin_clk_2_, bottom_width_0_height_0_subtile_15__pin_clk_3_, bottom_width_0_height_0_subtile_15__pin_clk_4_, bottom_width_0_height_0_subtile_15__pin_clk_5_, bottom_width_0_height_0_subtile_15__pin_clk_6_, bottom_width_0_height_0_subtile_15__pin_clk_7_, bottom_width_0_height_0_subtile_15__pin_clk_8_, bottom_width_0_height_0_subtile_15__pin_clk_9_, bottom_width_0_height_0_subtile_15__pin_clk_10_, bottom_width_0_height_0_subtile_15__pin_clk_11_, bottom_width_0_height_0_subtile_15__pin_clk_12_, bottom_width_0_height_0_subtile_15__pin_clk_13_, bottom_width_0_height_0_subtile_15__pin_clk_14_, bottom_width_0_height_0_subtile_15__pin_clk_15_}),
		.ccff_head(logical_tile_io_corner_mode_io_corner__14_ccff_tail),
		.io_corner_a2f_o({right_width_0_height_0_subtile_15__pin_a2f_o_0_, right_width_0_height_0_subtile_15__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_15__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_corner_mode_io_corner__15_ccff_tail));

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__16 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[16]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[16]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[16]),
		.io_corner_f2a_i(top_width_0_height_0_subtile_16__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_16__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_16__pin_clk_0_, bottom_width_0_height_0_subtile_16__pin_clk_1_, bottom_width_0_height_0_subtile_16__pin_clk_2_, bottom_width_0_height_0_subtile_16__pin_clk_3_, bottom_width_0_height_0_subtile_16__pin_clk_4_, bottom_width_0_height_0_subtile_16__pin_clk_5_, bottom_width_0_height_0_subtile_16__pin_clk_6_, bottom_width_0_height_0_subtile_16__pin_clk_7_, bottom_width_0_height_0_subtile_16__pin_clk_8_, bottom_width_0_height_0_subtile_16__pin_clk_9_, bottom_width_0_height_0_subtile_16__pin_clk_10_, bottom_width_0_height_0_subtile_16__pin_clk_11_, bottom_width_0_height_0_subtile_16__pin_clk_12_, bottom_width_0_height_0_subtile_16__pin_clk_13_, bottom_width_0_height_0_subtile_16__pin_clk_14_, bottom_width_0_height_0_subtile_16__pin_clk_15_}),
		.ccff_head(logical_tile_io_corner_mode_io_corner__15_ccff_tail),
		.io_corner_a2f_o({right_width_0_height_0_subtile_16__pin_a2f_o_0_, right_width_0_height_0_subtile_16__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_16__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_corner_mode_io_corner__16_ccff_tail));

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__17 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[17]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[17]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[17]),
		.io_corner_f2a_i(top_width_0_height_0_subtile_17__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_17__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_17__pin_clk_0_, bottom_width_0_height_0_subtile_17__pin_clk_1_, bottom_width_0_height_0_subtile_17__pin_clk_2_, bottom_width_0_height_0_subtile_17__pin_clk_3_, bottom_width_0_height_0_subtile_17__pin_clk_4_, bottom_width_0_height_0_subtile_17__pin_clk_5_, bottom_width_0_height_0_subtile_17__pin_clk_6_, bottom_width_0_height_0_subtile_17__pin_clk_7_, bottom_width_0_height_0_subtile_17__pin_clk_8_, bottom_width_0_height_0_subtile_17__pin_clk_9_, bottom_width_0_height_0_subtile_17__pin_clk_10_, bottom_width_0_height_0_subtile_17__pin_clk_11_, bottom_width_0_height_0_subtile_17__pin_clk_12_, bottom_width_0_height_0_subtile_17__pin_clk_13_, bottom_width_0_height_0_subtile_17__pin_clk_14_, bottom_width_0_height_0_subtile_17__pin_clk_15_}),
		.ccff_head(logical_tile_io_corner_mode_io_corner__16_ccff_tail),
		.io_corner_a2f_o({right_width_0_height_0_subtile_17__pin_a2f_o_0_, right_width_0_height_0_subtile_17__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_17__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_corner_mode_io_corner__17_ccff_tail));

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__18 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[18]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[18]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[18]),
		.io_corner_f2a_i(top_width_0_height_0_subtile_18__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_18__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_18__pin_clk_0_, bottom_width_0_height_0_subtile_18__pin_clk_1_, bottom_width_0_height_0_subtile_18__pin_clk_2_, bottom_width_0_height_0_subtile_18__pin_clk_3_, bottom_width_0_height_0_subtile_18__pin_clk_4_, bottom_width_0_height_0_subtile_18__pin_clk_5_, bottom_width_0_height_0_subtile_18__pin_clk_6_, bottom_width_0_height_0_subtile_18__pin_clk_7_, bottom_width_0_height_0_subtile_18__pin_clk_8_, bottom_width_0_height_0_subtile_18__pin_clk_9_, bottom_width_0_height_0_subtile_18__pin_clk_10_, bottom_width_0_height_0_subtile_18__pin_clk_11_, bottom_width_0_height_0_subtile_18__pin_clk_12_, bottom_width_0_height_0_subtile_18__pin_clk_13_, bottom_width_0_height_0_subtile_18__pin_clk_14_, bottom_width_0_height_0_subtile_18__pin_clk_15_}),
		.ccff_head(logical_tile_io_corner_mode_io_corner__17_ccff_tail),
		.io_corner_a2f_o({right_width_0_height_0_subtile_18__pin_a2f_o_0_, right_width_0_height_0_subtile_18__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_18__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_corner_mode_io_corner__18_ccff_tail));

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__19 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[19]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[19]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[19]),
		.io_corner_f2a_i(top_width_0_height_0_subtile_19__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_19__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_19__pin_clk_0_, bottom_width_0_height_0_subtile_19__pin_clk_1_, bottom_width_0_height_0_subtile_19__pin_clk_2_, bottom_width_0_height_0_subtile_19__pin_clk_3_, bottom_width_0_height_0_subtile_19__pin_clk_4_, bottom_width_0_height_0_subtile_19__pin_clk_5_, bottom_width_0_height_0_subtile_19__pin_clk_6_, bottom_width_0_height_0_subtile_19__pin_clk_7_, bottom_width_0_height_0_subtile_19__pin_clk_8_, bottom_width_0_height_0_subtile_19__pin_clk_9_, bottom_width_0_height_0_subtile_19__pin_clk_10_, bottom_width_0_height_0_subtile_19__pin_clk_11_, bottom_width_0_height_0_subtile_19__pin_clk_12_, bottom_width_0_height_0_subtile_19__pin_clk_13_, bottom_width_0_height_0_subtile_19__pin_clk_14_, bottom_width_0_height_0_subtile_19__pin_clk_15_}),
		.ccff_head(logical_tile_io_corner_mode_io_corner__18_ccff_tail),
		.io_corner_a2f_o({right_width_0_height_0_subtile_19__pin_a2f_o_0_, right_width_0_height_0_subtile_19__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_19__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_corner_mode_io_corner__19_ccff_tail));

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__20 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[20]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[20]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[20]),
		.io_corner_f2a_i(top_width_0_height_0_subtile_20__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_20__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_20__pin_clk_0_, bottom_width_0_height_0_subtile_20__pin_clk_1_, bottom_width_0_height_0_subtile_20__pin_clk_2_, bottom_width_0_height_0_subtile_20__pin_clk_3_, bottom_width_0_height_0_subtile_20__pin_clk_4_, bottom_width_0_height_0_subtile_20__pin_clk_5_, bottom_width_0_height_0_subtile_20__pin_clk_6_, bottom_width_0_height_0_subtile_20__pin_clk_7_, bottom_width_0_height_0_subtile_20__pin_clk_8_, bottom_width_0_height_0_subtile_20__pin_clk_9_, bottom_width_0_height_0_subtile_20__pin_clk_10_, bottom_width_0_height_0_subtile_20__pin_clk_11_, bottom_width_0_height_0_subtile_20__pin_clk_12_, bottom_width_0_height_0_subtile_20__pin_clk_13_, bottom_width_0_height_0_subtile_20__pin_clk_14_, bottom_width_0_height_0_subtile_20__pin_clk_15_}),
		.ccff_head(logical_tile_io_corner_mode_io_corner__19_ccff_tail),
		.io_corner_a2f_o({right_width_0_height_0_subtile_20__pin_a2f_o_0_, right_width_0_height_0_subtile_20__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_20__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_corner_mode_io_corner__20_ccff_tail));

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__21 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[21]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[21]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[21]),
		.io_corner_f2a_i(top_width_0_height_0_subtile_21__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_21__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_21__pin_clk_0_, bottom_width_0_height_0_subtile_21__pin_clk_1_, bottom_width_0_height_0_subtile_21__pin_clk_2_, bottom_width_0_height_0_subtile_21__pin_clk_3_, bottom_width_0_height_0_subtile_21__pin_clk_4_, bottom_width_0_height_0_subtile_21__pin_clk_5_, bottom_width_0_height_0_subtile_21__pin_clk_6_, bottom_width_0_height_0_subtile_21__pin_clk_7_, bottom_width_0_height_0_subtile_21__pin_clk_8_, bottom_width_0_height_0_subtile_21__pin_clk_9_, bottom_width_0_height_0_subtile_21__pin_clk_10_, bottom_width_0_height_0_subtile_21__pin_clk_11_, bottom_width_0_height_0_subtile_21__pin_clk_12_, bottom_width_0_height_0_subtile_21__pin_clk_13_, bottom_width_0_height_0_subtile_21__pin_clk_14_, bottom_width_0_height_0_subtile_21__pin_clk_15_}),
		.ccff_head(logical_tile_io_corner_mode_io_corner__20_ccff_tail),
		.io_corner_a2f_o({right_width_0_height_0_subtile_21__pin_a2f_o_0_, right_width_0_height_0_subtile_21__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_21__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_corner_mode_io_corner__21_ccff_tail));

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__22 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[22]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[22]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[22]),
		.io_corner_f2a_i(top_width_0_height_0_subtile_22__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_22__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_22__pin_clk_0_, bottom_width_0_height_0_subtile_22__pin_clk_1_, bottom_width_0_height_0_subtile_22__pin_clk_2_, bottom_width_0_height_0_subtile_22__pin_clk_3_, bottom_width_0_height_0_subtile_22__pin_clk_4_, bottom_width_0_height_0_subtile_22__pin_clk_5_, bottom_width_0_height_0_subtile_22__pin_clk_6_, bottom_width_0_height_0_subtile_22__pin_clk_7_, bottom_width_0_height_0_subtile_22__pin_clk_8_, bottom_width_0_height_0_subtile_22__pin_clk_9_, bottom_width_0_height_0_subtile_22__pin_clk_10_, bottom_width_0_height_0_subtile_22__pin_clk_11_, bottom_width_0_height_0_subtile_22__pin_clk_12_, bottom_width_0_height_0_subtile_22__pin_clk_13_, bottom_width_0_height_0_subtile_22__pin_clk_14_, bottom_width_0_height_0_subtile_22__pin_clk_15_}),
		.ccff_head(logical_tile_io_corner_mode_io_corner__21_ccff_tail),
		.io_corner_a2f_o({right_width_0_height_0_subtile_22__pin_a2f_o_0_, right_width_0_height_0_subtile_22__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_22__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_corner_mode_io_corner__22_ccff_tail));

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__23 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[23]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[23]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[23]),
		.io_corner_f2a_i(top_width_0_height_0_subtile_23__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_23__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_23__pin_clk_0_, bottom_width_0_height_0_subtile_23__pin_clk_1_, bottom_width_0_height_0_subtile_23__pin_clk_2_, bottom_width_0_height_0_subtile_23__pin_clk_3_, bottom_width_0_height_0_subtile_23__pin_clk_4_, bottom_width_0_height_0_subtile_23__pin_clk_5_, bottom_width_0_height_0_subtile_23__pin_clk_6_, bottom_width_0_height_0_subtile_23__pin_clk_7_, bottom_width_0_height_0_subtile_23__pin_clk_8_, bottom_width_0_height_0_subtile_23__pin_clk_9_, bottom_width_0_height_0_subtile_23__pin_clk_10_, bottom_width_0_height_0_subtile_23__pin_clk_11_, bottom_width_0_height_0_subtile_23__pin_clk_12_, bottom_width_0_height_0_subtile_23__pin_clk_13_, bottom_width_0_height_0_subtile_23__pin_clk_14_, bottom_width_0_height_0_subtile_23__pin_clk_15_}),
		.ccff_head(logical_tile_io_corner_mode_io_corner__22_ccff_tail),
		.io_corner_a2f_o({right_width_0_height_0_subtile_23__pin_a2f_o_0_, right_width_0_height_0_subtile_23__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_23__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_corner_mode_io_corner__23_ccff_tail));

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__24 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[24]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[24]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[24]),
		.io_corner_f2a_i(top_width_0_height_0_subtile_24__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_24__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_24__pin_clk_0_, bottom_width_0_height_0_subtile_24__pin_clk_1_, bottom_width_0_height_0_subtile_24__pin_clk_2_, bottom_width_0_height_0_subtile_24__pin_clk_3_, bottom_width_0_height_0_subtile_24__pin_clk_4_, bottom_width_0_height_0_subtile_24__pin_clk_5_, bottom_width_0_height_0_subtile_24__pin_clk_6_, bottom_width_0_height_0_subtile_24__pin_clk_7_, bottom_width_0_height_0_subtile_24__pin_clk_8_, bottom_width_0_height_0_subtile_24__pin_clk_9_, bottom_width_0_height_0_subtile_24__pin_clk_10_, bottom_width_0_height_0_subtile_24__pin_clk_11_, bottom_width_0_height_0_subtile_24__pin_clk_12_, bottom_width_0_height_0_subtile_24__pin_clk_13_, bottom_width_0_height_0_subtile_24__pin_clk_14_, bottom_width_0_height_0_subtile_24__pin_clk_15_}),
		.ccff_head(logical_tile_io_corner_mode_io_corner__23_ccff_tail),
		.io_corner_a2f_o({right_width_0_height_0_subtile_24__pin_a2f_o_0_, right_width_0_height_0_subtile_24__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_24__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_corner_mode_io_corner__24_ccff_tail));

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__25 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[25]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[25]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[25]),
		.io_corner_f2a_i(top_width_0_height_0_subtile_25__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_25__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_25__pin_clk_0_, bottom_width_0_height_0_subtile_25__pin_clk_1_, bottom_width_0_height_0_subtile_25__pin_clk_2_, bottom_width_0_height_0_subtile_25__pin_clk_3_, bottom_width_0_height_0_subtile_25__pin_clk_4_, bottom_width_0_height_0_subtile_25__pin_clk_5_, bottom_width_0_height_0_subtile_25__pin_clk_6_, bottom_width_0_height_0_subtile_25__pin_clk_7_, bottom_width_0_height_0_subtile_25__pin_clk_8_, bottom_width_0_height_0_subtile_25__pin_clk_9_, bottom_width_0_height_0_subtile_25__pin_clk_10_, bottom_width_0_height_0_subtile_25__pin_clk_11_, bottom_width_0_height_0_subtile_25__pin_clk_12_, bottom_width_0_height_0_subtile_25__pin_clk_13_, bottom_width_0_height_0_subtile_25__pin_clk_14_, bottom_width_0_height_0_subtile_25__pin_clk_15_}),
		.ccff_head(logical_tile_io_corner_mode_io_corner__24_ccff_tail),
		.io_corner_a2f_o({right_width_0_height_0_subtile_25__pin_a2f_o_0_, right_width_0_height_0_subtile_25__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_25__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_corner_mode_io_corner__25_ccff_tail));

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__26 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[26]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[26]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[26]),
		.io_corner_f2a_i(top_width_0_height_0_subtile_26__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_26__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_26__pin_clk_0_, bottom_width_0_height_0_subtile_26__pin_clk_1_, bottom_width_0_height_0_subtile_26__pin_clk_2_, bottom_width_0_height_0_subtile_26__pin_clk_3_, bottom_width_0_height_0_subtile_26__pin_clk_4_, bottom_width_0_height_0_subtile_26__pin_clk_5_, bottom_width_0_height_0_subtile_26__pin_clk_6_, bottom_width_0_height_0_subtile_26__pin_clk_7_, bottom_width_0_height_0_subtile_26__pin_clk_8_, bottom_width_0_height_0_subtile_26__pin_clk_9_, bottom_width_0_height_0_subtile_26__pin_clk_10_, bottom_width_0_height_0_subtile_26__pin_clk_11_, bottom_width_0_height_0_subtile_26__pin_clk_12_, bottom_width_0_height_0_subtile_26__pin_clk_13_, bottom_width_0_height_0_subtile_26__pin_clk_14_, bottom_width_0_height_0_subtile_26__pin_clk_15_}),
		.ccff_head(logical_tile_io_corner_mode_io_corner__25_ccff_tail),
		.io_corner_a2f_o({right_width_0_height_0_subtile_26__pin_a2f_o_0_, right_width_0_height_0_subtile_26__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_26__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_corner_mode_io_corner__26_ccff_tail));

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__27 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[27]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[27]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[27]),
		.io_corner_f2a_i(top_width_0_height_0_subtile_27__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_27__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_27__pin_clk_0_, bottom_width_0_height_0_subtile_27__pin_clk_1_, bottom_width_0_height_0_subtile_27__pin_clk_2_, bottom_width_0_height_0_subtile_27__pin_clk_3_, bottom_width_0_height_0_subtile_27__pin_clk_4_, bottom_width_0_height_0_subtile_27__pin_clk_5_, bottom_width_0_height_0_subtile_27__pin_clk_6_, bottom_width_0_height_0_subtile_27__pin_clk_7_, bottom_width_0_height_0_subtile_27__pin_clk_8_, bottom_width_0_height_0_subtile_27__pin_clk_9_, bottom_width_0_height_0_subtile_27__pin_clk_10_, bottom_width_0_height_0_subtile_27__pin_clk_11_, bottom_width_0_height_0_subtile_27__pin_clk_12_, bottom_width_0_height_0_subtile_27__pin_clk_13_, bottom_width_0_height_0_subtile_27__pin_clk_14_, bottom_width_0_height_0_subtile_27__pin_clk_15_}),
		.ccff_head(logical_tile_io_corner_mode_io_corner__26_ccff_tail),
		.io_corner_a2f_o({right_width_0_height_0_subtile_27__pin_a2f_o_0_, right_width_0_height_0_subtile_27__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_27__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_corner_mode_io_corner__27_ccff_tail));

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__28 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[28]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[28]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[28]),
		.io_corner_f2a_i(top_width_0_height_0_subtile_28__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_28__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_28__pin_clk_0_, bottom_width_0_height_0_subtile_28__pin_clk_1_, bottom_width_0_height_0_subtile_28__pin_clk_2_, bottom_width_0_height_0_subtile_28__pin_clk_3_, bottom_width_0_height_0_subtile_28__pin_clk_4_, bottom_width_0_height_0_subtile_28__pin_clk_5_, bottom_width_0_height_0_subtile_28__pin_clk_6_, bottom_width_0_height_0_subtile_28__pin_clk_7_, bottom_width_0_height_0_subtile_28__pin_clk_8_, bottom_width_0_height_0_subtile_28__pin_clk_9_, bottom_width_0_height_0_subtile_28__pin_clk_10_, bottom_width_0_height_0_subtile_28__pin_clk_11_, bottom_width_0_height_0_subtile_28__pin_clk_12_, bottom_width_0_height_0_subtile_28__pin_clk_13_, bottom_width_0_height_0_subtile_28__pin_clk_14_, bottom_width_0_height_0_subtile_28__pin_clk_15_}),
		.ccff_head(logical_tile_io_corner_mode_io_corner__27_ccff_tail),
		.io_corner_a2f_o({right_width_0_height_0_subtile_28__pin_a2f_o_0_, right_width_0_height_0_subtile_28__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_28__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_corner_mode_io_corner__28_ccff_tail));

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__29 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[29]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[29]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[29]),
		.io_corner_f2a_i(top_width_0_height_0_subtile_29__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_29__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_29__pin_clk_0_, bottom_width_0_height_0_subtile_29__pin_clk_1_, bottom_width_0_height_0_subtile_29__pin_clk_2_, bottom_width_0_height_0_subtile_29__pin_clk_3_, bottom_width_0_height_0_subtile_29__pin_clk_4_, bottom_width_0_height_0_subtile_29__pin_clk_5_, bottom_width_0_height_0_subtile_29__pin_clk_6_, bottom_width_0_height_0_subtile_29__pin_clk_7_, bottom_width_0_height_0_subtile_29__pin_clk_8_, bottom_width_0_height_0_subtile_29__pin_clk_9_, bottom_width_0_height_0_subtile_29__pin_clk_10_, bottom_width_0_height_0_subtile_29__pin_clk_11_, bottom_width_0_height_0_subtile_29__pin_clk_12_, bottom_width_0_height_0_subtile_29__pin_clk_13_, bottom_width_0_height_0_subtile_29__pin_clk_14_, bottom_width_0_height_0_subtile_29__pin_clk_15_}),
		.ccff_head(logical_tile_io_corner_mode_io_corner__28_ccff_tail),
		.io_corner_a2f_o({right_width_0_height_0_subtile_29__pin_a2f_o_0_, right_width_0_height_0_subtile_29__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_29__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_corner_mode_io_corner__29_ccff_tail));

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__30 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[30]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[30]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[30]),
		.io_corner_f2a_i(top_width_0_height_0_subtile_30__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_30__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_30__pin_clk_0_, bottom_width_0_height_0_subtile_30__pin_clk_1_, bottom_width_0_height_0_subtile_30__pin_clk_2_, bottom_width_0_height_0_subtile_30__pin_clk_3_, bottom_width_0_height_0_subtile_30__pin_clk_4_, bottom_width_0_height_0_subtile_30__pin_clk_5_, bottom_width_0_height_0_subtile_30__pin_clk_6_, bottom_width_0_height_0_subtile_30__pin_clk_7_, bottom_width_0_height_0_subtile_30__pin_clk_8_, bottom_width_0_height_0_subtile_30__pin_clk_9_, bottom_width_0_height_0_subtile_30__pin_clk_10_, bottom_width_0_height_0_subtile_30__pin_clk_11_, bottom_width_0_height_0_subtile_30__pin_clk_12_, bottom_width_0_height_0_subtile_30__pin_clk_13_, bottom_width_0_height_0_subtile_30__pin_clk_14_, bottom_width_0_height_0_subtile_30__pin_clk_15_}),
		.ccff_head(logical_tile_io_corner_mode_io_corner__29_ccff_tail),
		.io_corner_a2f_o({top_width_0_height_0_subtile_30__pin_a2f_o_0_, top_width_0_height_0_subtile_30__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_30__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_corner_mode_io_corner__30_ccff_tail));

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__31 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[31]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[31]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[31]),
		.io_corner_f2a_i(top_width_0_height_0_subtile_31__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_31__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_31__pin_clk_0_, bottom_width_0_height_0_subtile_31__pin_clk_1_, bottom_width_0_height_0_subtile_31__pin_clk_2_, bottom_width_0_height_0_subtile_31__pin_clk_3_, bottom_width_0_height_0_subtile_31__pin_clk_4_, bottom_width_0_height_0_subtile_31__pin_clk_5_, bottom_width_0_height_0_subtile_31__pin_clk_6_, bottom_width_0_height_0_subtile_31__pin_clk_7_, bottom_width_0_height_0_subtile_31__pin_clk_8_, bottom_width_0_height_0_subtile_31__pin_clk_9_, bottom_width_0_height_0_subtile_31__pin_clk_10_, bottom_width_0_height_0_subtile_31__pin_clk_11_, bottom_width_0_height_0_subtile_31__pin_clk_12_, bottom_width_0_height_0_subtile_31__pin_clk_13_, bottom_width_0_height_0_subtile_31__pin_clk_14_, bottom_width_0_height_0_subtile_31__pin_clk_15_}),
		.ccff_head(logical_tile_io_corner_mode_io_corner__30_ccff_tail),
		.io_corner_a2f_o({top_width_0_height_0_subtile_31__pin_a2f_o_0_, top_width_0_height_0_subtile_31__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_31__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_corner_mode_io_corner__31_ccff_tail));

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__32 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[32]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[32]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[32]),
		.io_corner_f2a_i(top_width_0_height_0_subtile_32__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_32__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_32__pin_clk_0_, bottom_width_0_height_0_subtile_32__pin_clk_1_, bottom_width_0_height_0_subtile_32__pin_clk_2_, bottom_width_0_height_0_subtile_32__pin_clk_3_, bottom_width_0_height_0_subtile_32__pin_clk_4_, bottom_width_0_height_0_subtile_32__pin_clk_5_, bottom_width_0_height_0_subtile_32__pin_clk_6_, bottom_width_0_height_0_subtile_32__pin_clk_7_, bottom_width_0_height_0_subtile_32__pin_clk_8_, bottom_width_0_height_0_subtile_32__pin_clk_9_, bottom_width_0_height_0_subtile_32__pin_clk_10_, bottom_width_0_height_0_subtile_32__pin_clk_11_, bottom_width_0_height_0_subtile_32__pin_clk_12_, bottom_width_0_height_0_subtile_32__pin_clk_13_, bottom_width_0_height_0_subtile_32__pin_clk_14_, bottom_width_0_height_0_subtile_32__pin_clk_15_}),
		.ccff_head(logical_tile_io_corner_mode_io_corner__31_ccff_tail),
		.io_corner_a2f_o({top_width_0_height_0_subtile_32__pin_a2f_o_0_, top_width_0_height_0_subtile_32__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_32__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_corner_mode_io_corner__32_ccff_tail));

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__33 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[33]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[33]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[33]),
		.io_corner_f2a_i(top_width_0_height_0_subtile_33__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_33__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_33__pin_clk_0_, bottom_width_0_height_0_subtile_33__pin_clk_1_, bottom_width_0_height_0_subtile_33__pin_clk_2_, bottom_width_0_height_0_subtile_33__pin_clk_3_, bottom_width_0_height_0_subtile_33__pin_clk_4_, bottom_width_0_height_0_subtile_33__pin_clk_5_, bottom_width_0_height_0_subtile_33__pin_clk_6_, bottom_width_0_height_0_subtile_33__pin_clk_7_, bottom_width_0_height_0_subtile_33__pin_clk_8_, bottom_width_0_height_0_subtile_33__pin_clk_9_, bottom_width_0_height_0_subtile_33__pin_clk_10_, bottom_width_0_height_0_subtile_33__pin_clk_11_, bottom_width_0_height_0_subtile_33__pin_clk_12_, bottom_width_0_height_0_subtile_33__pin_clk_13_, bottom_width_0_height_0_subtile_33__pin_clk_14_, bottom_width_0_height_0_subtile_33__pin_clk_15_}),
		.ccff_head(logical_tile_io_corner_mode_io_corner__32_ccff_tail),
		.io_corner_a2f_o({top_width_0_height_0_subtile_33__pin_a2f_o_0_, top_width_0_height_0_subtile_33__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_33__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_corner_mode_io_corner__33_ccff_tail));

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__34 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[34]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[34]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[34]),
		.io_corner_f2a_i(top_width_0_height_0_subtile_34__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_34__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_34__pin_clk_0_, bottom_width_0_height_0_subtile_34__pin_clk_1_, bottom_width_0_height_0_subtile_34__pin_clk_2_, bottom_width_0_height_0_subtile_34__pin_clk_3_, bottom_width_0_height_0_subtile_34__pin_clk_4_, bottom_width_0_height_0_subtile_34__pin_clk_5_, bottom_width_0_height_0_subtile_34__pin_clk_6_, bottom_width_0_height_0_subtile_34__pin_clk_7_, bottom_width_0_height_0_subtile_34__pin_clk_8_, bottom_width_0_height_0_subtile_34__pin_clk_9_, bottom_width_0_height_0_subtile_34__pin_clk_10_, bottom_width_0_height_0_subtile_34__pin_clk_11_, bottom_width_0_height_0_subtile_34__pin_clk_12_, bottom_width_0_height_0_subtile_34__pin_clk_13_, bottom_width_0_height_0_subtile_34__pin_clk_14_, bottom_width_0_height_0_subtile_34__pin_clk_15_}),
		.ccff_head(logical_tile_io_corner_mode_io_corner__33_ccff_tail),
		.io_corner_a2f_o({top_width_0_height_0_subtile_34__pin_a2f_o_0_, top_width_0_height_0_subtile_34__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_34__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_corner_mode_io_corner__34_ccff_tail));

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__35 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[35]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[35]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[35]),
		.io_corner_f2a_i(top_width_0_height_0_subtile_35__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_35__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_35__pin_clk_0_, bottom_width_0_height_0_subtile_35__pin_clk_1_, bottom_width_0_height_0_subtile_35__pin_clk_2_, bottom_width_0_height_0_subtile_35__pin_clk_3_, bottom_width_0_height_0_subtile_35__pin_clk_4_, bottom_width_0_height_0_subtile_35__pin_clk_5_, bottom_width_0_height_0_subtile_35__pin_clk_6_, bottom_width_0_height_0_subtile_35__pin_clk_7_, bottom_width_0_height_0_subtile_35__pin_clk_8_, bottom_width_0_height_0_subtile_35__pin_clk_9_, bottom_width_0_height_0_subtile_35__pin_clk_10_, bottom_width_0_height_0_subtile_35__pin_clk_11_, bottom_width_0_height_0_subtile_35__pin_clk_12_, bottom_width_0_height_0_subtile_35__pin_clk_13_, bottom_width_0_height_0_subtile_35__pin_clk_14_, bottom_width_0_height_0_subtile_35__pin_clk_15_}),
		.ccff_head(logical_tile_io_corner_mode_io_corner__34_ccff_tail),
		.io_corner_a2f_o({top_width_0_height_0_subtile_35__pin_a2f_o_0_, top_width_0_height_0_subtile_35__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_35__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_corner_mode_io_corner__35_ccff_tail));

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__36 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[36]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[36]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[36]),
		.io_corner_f2a_i(top_width_0_height_0_subtile_36__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_36__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_36__pin_clk_0_, bottom_width_0_height_0_subtile_36__pin_clk_1_, bottom_width_0_height_0_subtile_36__pin_clk_2_, bottom_width_0_height_0_subtile_36__pin_clk_3_, bottom_width_0_height_0_subtile_36__pin_clk_4_, bottom_width_0_height_0_subtile_36__pin_clk_5_, bottom_width_0_height_0_subtile_36__pin_clk_6_, bottom_width_0_height_0_subtile_36__pin_clk_7_, bottom_width_0_height_0_subtile_36__pin_clk_8_, bottom_width_0_height_0_subtile_36__pin_clk_9_, bottom_width_0_height_0_subtile_36__pin_clk_10_, bottom_width_0_height_0_subtile_36__pin_clk_11_, bottom_width_0_height_0_subtile_36__pin_clk_12_, bottom_width_0_height_0_subtile_36__pin_clk_13_, bottom_width_0_height_0_subtile_36__pin_clk_14_, bottom_width_0_height_0_subtile_36__pin_clk_15_}),
		.ccff_head(logical_tile_io_corner_mode_io_corner__35_ccff_tail),
		.io_corner_a2f_o({top_width_0_height_0_subtile_36__pin_a2f_o_0_, top_width_0_height_0_subtile_36__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_36__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_corner_mode_io_corner__36_ccff_tail));

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__37 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[37]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[37]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[37]),
		.io_corner_f2a_i(top_width_0_height_0_subtile_37__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_37__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_37__pin_clk_0_, bottom_width_0_height_0_subtile_37__pin_clk_1_, bottom_width_0_height_0_subtile_37__pin_clk_2_, bottom_width_0_height_0_subtile_37__pin_clk_3_, bottom_width_0_height_0_subtile_37__pin_clk_4_, bottom_width_0_height_0_subtile_37__pin_clk_5_, bottom_width_0_height_0_subtile_37__pin_clk_6_, bottom_width_0_height_0_subtile_37__pin_clk_7_, bottom_width_0_height_0_subtile_37__pin_clk_8_, bottom_width_0_height_0_subtile_37__pin_clk_9_, bottom_width_0_height_0_subtile_37__pin_clk_10_, bottom_width_0_height_0_subtile_37__pin_clk_11_, bottom_width_0_height_0_subtile_37__pin_clk_12_, bottom_width_0_height_0_subtile_37__pin_clk_13_, bottom_width_0_height_0_subtile_37__pin_clk_14_, bottom_width_0_height_0_subtile_37__pin_clk_15_}),
		.ccff_head(logical_tile_io_corner_mode_io_corner__36_ccff_tail),
		.io_corner_a2f_o({top_width_0_height_0_subtile_37__pin_a2f_o_0_, top_width_0_height_0_subtile_37__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_37__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_corner_mode_io_corner__37_ccff_tail));

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__38 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[38]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[38]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[38]),
		.io_corner_f2a_i(top_width_0_height_0_subtile_38__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_38__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_38__pin_clk_0_, bottom_width_0_height_0_subtile_38__pin_clk_1_, bottom_width_0_height_0_subtile_38__pin_clk_2_, bottom_width_0_height_0_subtile_38__pin_clk_3_, bottom_width_0_height_0_subtile_38__pin_clk_4_, bottom_width_0_height_0_subtile_38__pin_clk_5_, bottom_width_0_height_0_subtile_38__pin_clk_6_, bottom_width_0_height_0_subtile_38__pin_clk_7_, bottom_width_0_height_0_subtile_38__pin_clk_8_, bottom_width_0_height_0_subtile_38__pin_clk_9_, bottom_width_0_height_0_subtile_38__pin_clk_10_, bottom_width_0_height_0_subtile_38__pin_clk_11_, bottom_width_0_height_0_subtile_38__pin_clk_12_, bottom_width_0_height_0_subtile_38__pin_clk_13_, bottom_width_0_height_0_subtile_38__pin_clk_14_, bottom_width_0_height_0_subtile_38__pin_clk_15_}),
		.ccff_head(logical_tile_io_corner_mode_io_corner__37_ccff_tail),
		.io_corner_a2f_o({top_width_0_height_0_subtile_38__pin_a2f_o_0_, top_width_0_height_0_subtile_38__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_38__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_corner_mode_io_corner__38_ccff_tail));

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__39 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[39]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[39]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[39]),
		.io_corner_f2a_i(top_width_0_height_0_subtile_39__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_39__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_39__pin_clk_0_, bottom_width_0_height_0_subtile_39__pin_clk_1_, bottom_width_0_height_0_subtile_39__pin_clk_2_, bottom_width_0_height_0_subtile_39__pin_clk_3_, bottom_width_0_height_0_subtile_39__pin_clk_4_, bottom_width_0_height_0_subtile_39__pin_clk_5_, bottom_width_0_height_0_subtile_39__pin_clk_6_, bottom_width_0_height_0_subtile_39__pin_clk_7_, bottom_width_0_height_0_subtile_39__pin_clk_8_, bottom_width_0_height_0_subtile_39__pin_clk_9_, bottom_width_0_height_0_subtile_39__pin_clk_10_, bottom_width_0_height_0_subtile_39__pin_clk_11_, bottom_width_0_height_0_subtile_39__pin_clk_12_, bottom_width_0_height_0_subtile_39__pin_clk_13_, bottom_width_0_height_0_subtile_39__pin_clk_14_, bottom_width_0_height_0_subtile_39__pin_clk_15_}),
		.ccff_head(logical_tile_io_corner_mode_io_corner__38_ccff_tail),
		.io_corner_a2f_o({top_width_0_height_0_subtile_39__pin_a2f_o_0_, top_width_0_height_0_subtile_39__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_39__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_corner_mode_io_corner__39_ccff_tail));

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__40 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[40]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[40]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[40]),
		.io_corner_f2a_i(top_width_0_height_0_subtile_40__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_40__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_40__pin_clk_0_, bottom_width_0_height_0_subtile_40__pin_clk_1_, bottom_width_0_height_0_subtile_40__pin_clk_2_, bottom_width_0_height_0_subtile_40__pin_clk_3_, bottom_width_0_height_0_subtile_40__pin_clk_4_, bottom_width_0_height_0_subtile_40__pin_clk_5_, bottom_width_0_height_0_subtile_40__pin_clk_6_, bottom_width_0_height_0_subtile_40__pin_clk_7_, bottom_width_0_height_0_subtile_40__pin_clk_8_, bottom_width_0_height_0_subtile_40__pin_clk_9_, bottom_width_0_height_0_subtile_40__pin_clk_10_, bottom_width_0_height_0_subtile_40__pin_clk_11_, bottom_width_0_height_0_subtile_40__pin_clk_12_, bottom_width_0_height_0_subtile_40__pin_clk_13_, bottom_width_0_height_0_subtile_40__pin_clk_14_, bottom_width_0_height_0_subtile_40__pin_clk_15_}),
		.ccff_head(logical_tile_io_corner_mode_io_corner__39_ccff_tail),
		.io_corner_a2f_o({top_width_0_height_0_subtile_40__pin_a2f_o_0_, top_width_0_height_0_subtile_40__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_40__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_corner_mode_io_corner__40_ccff_tail));

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__41 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[41]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[41]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[41]),
		.io_corner_f2a_i(top_width_0_height_0_subtile_41__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_41__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_41__pin_clk_0_, bottom_width_0_height_0_subtile_41__pin_clk_1_, bottom_width_0_height_0_subtile_41__pin_clk_2_, bottom_width_0_height_0_subtile_41__pin_clk_3_, bottom_width_0_height_0_subtile_41__pin_clk_4_, bottom_width_0_height_0_subtile_41__pin_clk_5_, bottom_width_0_height_0_subtile_41__pin_clk_6_, bottom_width_0_height_0_subtile_41__pin_clk_7_, bottom_width_0_height_0_subtile_41__pin_clk_8_, bottom_width_0_height_0_subtile_41__pin_clk_9_, bottom_width_0_height_0_subtile_41__pin_clk_10_, bottom_width_0_height_0_subtile_41__pin_clk_11_, bottom_width_0_height_0_subtile_41__pin_clk_12_, bottom_width_0_height_0_subtile_41__pin_clk_13_, bottom_width_0_height_0_subtile_41__pin_clk_14_, bottom_width_0_height_0_subtile_41__pin_clk_15_}),
		.ccff_head(logical_tile_io_corner_mode_io_corner__40_ccff_tail),
		.io_corner_a2f_o({top_width_0_height_0_subtile_41__pin_a2f_o_0_, top_width_0_height_0_subtile_41__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_41__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_corner_mode_io_corner__41_ccff_tail));

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__42 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[42]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[42]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[42]),
		.io_corner_f2a_i(top_width_0_height_0_subtile_42__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_42__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_42__pin_clk_0_, bottom_width_0_height_0_subtile_42__pin_clk_1_, bottom_width_0_height_0_subtile_42__pin_clk_2_, bottom_width_0_height_0_subtile_42__pin_clk_3_, bottom_width_0_height_0_subtile_42__pin_clk_4_, bottom_width_0_height_0_subtile_42__pin_clk_5_, bottom_width_0_height_0_subtile_42__pin_clk_6_, bottom_width_0_height_0_subtile_42__pin_clk_7_, bottom_width_0_height_0_subtile_42__pin_clk_8_, bottom_width_0_height_0_subtile_42__pin_clk_9_, bottom_width_0_height_0_subtile_42__pin_clk_10_, bottom_width_0_height_0_subtile_42__pin_clk_11_, bottom_width_0_height_0_subtile_42__pin_clk_12_, bottom_width_0_height_0_subtile_42__pin_clk_13_, bottom_width_0_height_0_subtile_42__pin_clk_14_, bottom_width_0_height_0_subtile_42__pin_clk_15_}),
		.ccff_head(logical_tile_io_corner_mode_io_corner__41_ccff_tail),
		.io_corner_a2f_o({top_width_0_height_0_subtile_42__pin_a2f_o_0_, top_width_0_height_0_subtile_42__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_42__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_corner_mode_io_corner__42_ccff_tail));

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__43 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[43]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[43]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[43]),
		.io_corner_f2a_i(top_width_0_height_0_subtile_43__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_43__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_43__pin_clk_0_, bottom_width_0_height_0_subtile_43__pin_clk_1_, bottom_width_0_height_0_subtile_43__pin_clk_2_, bottom_width_0_height_0_subtile_43__pin_clk_3_, bottom_width_0_height_0_subtile_43__pin_clk_4_, bottom_width_0_height_0_subtile_43__pin_clk_5_, bottom_width_0_height_0_subtile_43__pin_clk_6_, bottom_width_0_height_0_subtile_43__pin_clk_7_, bottom_width_0_height_0_subtile_43__pin_clk_8_, bottom_width_0_height_0_subtile_43__pin_clk_9_, bottom_width_0_height_0_subtile_43__pin_clk_10_, bottom_width_0_height_0_subtile_43__pin_clk_11_, bottom_width_0_height_0_subtile_43__pin_clk_12_, bottom_width_0_height_0_subtile_43__pin_clk_13_, bottom_width_0_height_0_subtile_43__pin_clk_14_, bottom_width_0_height_0_subtile_43__pin_clk_15_}),
		.ccff_head(logical_tile_io_corner_mode_io_corner__42_ccff_tail),
		.io_corner_a2f_o({top_width_0_height_0_subtile_43__pin_a2f_o_0_, top_width_0_height_0_subtile_43__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_43__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_corner_mode_io_corner__43_ccff_tail));

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__44 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[44]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[44]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[44]),
		.io_corner_f2a_i(top_width_0_height_0_subtile_44__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_44__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_44__pin_clk_0_, bottom_width_0_height_0_subtile_44__pin_clk_1_, bottom_width_0_height_0_subtile_44__pin_clk_2_, bottom_width_0_height_0_subtile_44__pin_clk_3_, bottom_width_0_height_0_subtile_44__pin_clk_4_, bottom_width_0_height_0_subtile_44__pin_clk_5_, bottom_width_0_height_0_subtile_44__pin_clk_6_, bottom_width_0_height_0_subtile_44__pin_clk_7_, bottom_width_0_height_0_subtile_44__pin_clk_8_, bottom_width_0_height_0_subtile_44__pin_clk_9_, bottom_width_0_height_0_subtile_44__pin_clk_10_, bottom_width_0_height_0_subtile_44__pin_clk_11_, bottom_width_0_height_0_subtile_44__pin_clk_12_, bottom_width_0_height_0_subtile_44__pin_clk_13_, bottom_width_0_height_0_subtile_44__pin_clk_14_, bottom_width_0_height_0_subtile_44__pin_clk_15_}),
		.ccff_head(logical_tile_io_corner_mode_io_corner__43_ccff_tail),
		.io_corner_a2f_o({top_width_0_height_0_subtile_44__pin_a2f_o_0_, top_width_0_height_0_subtile_44__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_44__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_corner_mode_io_corner__44_ccff_tail));

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__45 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[45]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[45]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[45]),
		.io_corner_f2a_i(top_width_0_height_0_subtile_45__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_45__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_45__pin_clk_0_, bottom_width_0_height_0_subtile_45__pin_clk_1_, bottom_width_0_height_0_subtile_45__pin_clk_2_, bottom_width_0_height_0_subtile_45__pin_clk_3_, bottom_width_0_height_0_subtile_45__pin_clk_4_, bottom_width_0_height_0_subtile_45__pin_clk_5_, bottom_width_0_height_0_subtile_45__pin_clk_6_, bottom_width_0_height_0_subtile_45__pin_clk_7_, bottom_width_0_height_0_subtile_45__pin_clk_8_, bottom_width_0_height_0_subtile_45__pin_clk_9_, bottom_width_0_height_0_subtile_45__pin_clk_10_, bottom_width_0_height_0_subtile_45__pin_clk_11_, bottom_width_0_height_0_subtile_45__pin_clk_12_, bottom_width_0_height_0_subtile_45__pin_clk_13_, bottom_width_0_height_0_subtile_45__pin_clk_14_, bottom_width_0_height_0_subtile_45__pin_clk_15_}),
		.ccff_head(logical_tile_io_corner_mode_io_corner__44_ccff_tail),
		.io_corner_a2f_o({top_width_0_height_0_subtile_45__pin_a2f_o_0_, top_width_0_height_0_subtile_45__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_45__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_corner_mode_io_corner__45_ccff_tail));

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__46 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[46]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[46]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[46]),
		.io_corner_f2a_i(top_width_0_height_0_subtile_46__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_46__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_46__pin_clk_0_, bottom_width_0_height_0_subtile_46__pin_clk_1_, bottom_width_0_height_0_subtile_46__pin_clk_2_, bottom_width_0_height_0_subtile_46__pin_clk_3_, bottom_width_0_height_0_subtile_46__pin_clk_4_, bottom_width_0_height_0_subtile_46__pin_clk_5_, bottom_width_0_height_0_subtile_46__pin_clk_6_, bottom_width_0_height_0_subtile_46__pin_clk_7_, bottom_width_0_height_0_subtile_46__pin_clk_8_, bottom_width_0_height_0_subtile_46__pin_clk_9_, bottom_width_0_height_0_subtile_46__pin_clk_10_, bottom_width_0_height_0_subtile_46__pin_clk_11_, bottom_width_0_height_0_subtile_46__pin_clk_12_, bottom_width_0_height_0_subtile_46__pin_clk_13_, bottom_width_0_height_0_subtile_46__pin_clk_14_, bottom_width_0_height_0_subtile_46__pin_clk_15_}),
		.ccff_head(logical_tile_io_corner_mode_io_corner__45_ccff_tail),
		.io_corner_a2f_o({top_width_0_height_0_subtile_46__pin_a2f_o_0_, top_width_0_height_0_subtile_46__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_46__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_corner_mode_io_corner__46_ccff_tail));

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__47 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[47]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[47]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[47]),
		.io_corner_f2a_i(top_width_0_height_0_subtile_47__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_47__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_47__pin_clk_0_, bottom_width_0_height_0_subtile_47__pin_clk_1_, bottom_width_0_height_0_subtile_47__pin_clk_2_, bottom_width_0_height_0_subtile_47__pin_clk_3_, bottom_width_0_height_0_subtile_47__pin_clk_4_, bottom_width_0_height_0_subtile_47__pin_clk_5_, bottom_width_0_height_0_subtile_47__pin_clk_6_, bottom_width_0_height_0_subtile_47__pin_clk_7_, bottom_width_0_height_0_subtile_47__pin_clk_8_, bottom_width_0_height_0_subtile_47__pin_clk_9_, bottom_width_0_height_0_subtile_47__pin_clk_10_, bottom_width_0_height_0_subtile_47__pin_clk_11_, bottom_width_0_height_0_subtile_47__pin_clk_12_, bottom_width_0_height_0_subtile_47__pin_clk_13_, bottom_width_0_height_0_subtile_47__pin_clk_14_, bottom_width_0_height_0_subtile_47__pin_clk_15_}),
		.ccff_head(logical_tile_io_corner_mode_io_corner__46_ccff_tail),
		.io_corner_a2f_o({top_width_0_height_0_subtile_47__pin_a2f_o_0_, top_width_0_height_0_subtile_47__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_47__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_corner_mode_io_corner__47_ccff_tail));

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__48 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[48]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[48]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[48]),
		.io_corner_f2a_i(top_width_0_height_0_subtile_48__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_48__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_48__pin_clk_0_, bottom_width_0_height_0_subtile_48__pin_clk_1_, bottom_width_0_height_0_subtile_48__pin_clk_2_, bottom_width_0_height_0_subtile_48__pin_clk_3_, bottom_width_0_height_0_subtile_48__pin_clk_4_, bottom_width_0_height_0_subtile_48__pin_clk_5_, bottom_width_0_height_0_subtile_48__pin_clk_6_, bottom_width_0_height_0_subtile_48__pin_clk_7_, bottom_width_0_height_0_subtile_48__pin_clk_8_, bottom_width_0_height_0_subtile_48__pin_clk_9_, bottom_width_0_height_0_subtile_48__pin_clk_10_, bottom_width_0_height_0_subtile_48__pin_clk_11_, bottom_width_0_height_0_subtile_48__pin_clk_12_, bottom_width_0_height_0_subtile_48__pin_clk_13_, bottom_width_0_height_0_subtile_48__pin_clk_14_, bottom_width_0_height_0_subtile_48__pin_clk_15_}),
		.ccff_head(logical_tile_io_corner_mode_io_corner__47_ccff_tail),
		.io_corner_a2f_o({top_width_0_height_0_subtile_48__pin_a2f_o_0_, top_width_0_height_0_subtile_48__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_48__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_corner_mode_io_corner__48_ccff_tail));

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__49 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[49]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[49]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[49]),
		.io_corner_f2a_i(top_width_0_height_0_subtile_49__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_49__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_49__pin_clk_0_, bottom_width_0_height_0_subtile_49__pin_clk_1_, bottom_width_0_height_0_subtile_49__pin_clk_2_, bottom_width_0_height_0_subtile_49__pin_clk_3_, bottom_width_0_height_0_subtile_49__pin_clk_4_, bottom_width_0_height_0_subtile_49__pin_clk_5_, bottom_width_0_height_0_subtile_49__pin_clk_6_, bottom_width_0_height_0_subtile_49__pin_clk_7_, bottom_width_0_height_0_subtile_49__pin_clk_8_, bottom_width_0_height_0_subtile_49__pin_clk_9_, bottom_width_0_height_0_subtile_49__pin_clk_10_, bottom_width_0_height_0_subtile_49__pin_clk_11_, bottom_width_0_height_0_subtile_49__pin_clk_12_, bottom_width_0_height_0_subtile_49__pin_clk_13_, bottom_width_0_height_0_subtile_49__pin_clk_14_, bottom_width_0_height_0_subtile_49__pin_clk_15_}),
		.ccff_head(logical_tile_io_corner_mode_io_corner__48_ccff_tail),
		.io_corner_a2f_o({top_width_0_height_0_subtile_49__pin_a2f_o_0_, top_width_0_height_0_subtile_49__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_49__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_corner_mode_io_corner__49_ccff_tail));

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__50 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[50]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[50]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[50]),
		.io_corner_f2a_i(top_width_0_height_0_subtile_50__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_50__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_50__pin_clk_0_, bottom_width_0_height_0_subtile_50__pin_clk_1_, bottom_width_0_height_0_subtile_50__pin_clk_2_, bottom_width_0_height_0_subtile_50__pin_clk_3_, bottom_width_0_height_0_subtile_50__pin_clk_4_, bottom_width_0_height_0_subtile_50__pin_clk_5_, bottom_width_0_height_0_subtile_50__pin_clk_6_, bottom_width_0_height_0_subtile_50__pin_clk_7_, bottom_width_0_height_0_subtile_50__pin_clk_8_, bottom_width_0_height_0_subtile_50__pin_clk_9_, bottom_width_0_height_0_subtile_50__pin_clk_10_, bottom_width_0_height_0_subtile_50__pin_clk_11_, bottom_width_0_height_0_subtile_50__pin_clk_12_, bottom_width_0_height_0_subtile_50__pin_clk_13_, bottom_width_0_height_0_subtile_50__pin_clk_14_, bottom_width_0_height_0_subtile_50__pin_clk_15_}),
		.ccff_head(logical_tile_io_corner_mode_io_corner__49_ccff_tail),
		.io_corner_a2f_o({top_width_0_height_0_subtile_50__pin_a2f_o_0_, top_width_0_height_0_subtile_50__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_50__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_corner_mode_io_corner__50_ccff_tail));

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__51 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[51]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[51]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[51]),
		.io_corner_f2a_i(top_width_0_height_0_subtile_51__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_51__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_51__pin_clk_0_, bottom_width_0_height_0_subtile_51__pin_clk_1_, bottom_width_0_height_0_subtile_51__pin_clk_2_, bottom_width_0_height_0_subtile_51__pin_clk_3_, bottom_width_0_height_0_subtile_51__pin_clk_4_, bottom_width_0_height_0_subtile_51__pin_clk_5_, bottom_width_0_height_0_subtile_51__pin_clk_6_, bottom_width_0_height_0_subtile_51__pin_clk_7_, bottom_width_0_height_0_subtile_51__pin_clk_8_, bottom_width_0_height_0_subtile_51__pin_clk_9_, bottom_width_0_height_0_subtile_51__pin_clk_10_, bottom_width_0_height_0_subtile_51__pin_clk_11_, bottom_width_0_height_0_subtile_51__pin_clk_12_, bottom_width_0_height_0_subtile_51__pin_clk_13_, bottom_width_0_height_0_subtile_51__pin_clk_14_, bottom_width_0_height_0_subtile_51__pin_clk_15_}),
		.ccff_head(logical_tile_io_corner_mode_io_corner__50_ccff_tail),
		.io_corner_a2f_o({top_width_0_height_0_subtile_51__pin_a2f_o_0_, top_width_0_height_0_subtile_51__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_51__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_corner_mode_io_corner__51_ccff_tail));

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__52 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[52]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[52]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[52]),
		.io_corner_f2a_i(top_width_0_height_0_subtile_52__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_52__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_52__pin_clk_0_, bottom_width_0_height_0_subtile_52__pin_clk_1_, bottom_width_0_height_0_subtile_52__pin_clk_2_, bottom_width_0_height_0_subtile_52__pin_clk_3_, bottom_width_0_height_0_subtile_52__pin_clk_4_, bottom_width_0_height_0_subtile_52__pin_clk_5_, bottom_width_0_height_0_subtile_52__pin_clk_6_, bottom_width_0_height_0_subtile_52__pin_clk_7_, bottom_width_0_height_0_subtile_52__pin_clk_8_, bottom_width_0_height_0_subtile_52__pin_clk_9_, bottom_width_0_height_0_subtile_52__pin_clk_10_, bottom_width_0_height_0_subtile_52__pin_clk_11_, bottom_width_0_height_0_subtile_52__pin_clk_12_, bottom_width_0_height_0_subtile_52__pin_clk_13_, bottom_width_0_height_0_subtile_52__pin_clk_14_, bottom_width_0_height_0_subtile_52__pin_clk_15_}),
		.ccff_head(logical_tile_io_corner_mode_io_corner__51_ccff_tail),
		.io_corner_a2f_o({top_width_0_height_0_subtile_52__pin_a2f_o_0_, top_width_0_height_0_subtile_52__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_52__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_corner_mode_io_corner__52_ccff_tail));

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__53 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[53]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[53]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[53]),
		.io_corner_f2a_i(top_width_0_height_0_subtile_53__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_53__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_53__pin_clk_0_, bottom_width_0_height_0_subtile_53__pin_clk_1_, bottom_width_0_height_0_subtile_53__pin_clk_2_, bottom_width_0_height_0_subtile_53__pin_clk_3_, bottom_width_0_height_0_subtile_53__pin_clk_4_, bottom_width_0_height_0_subtile_53__pin_clk_5_, bottom_width_0_height_0_subtile_53__pin_clk_6_, bottom_width_0_height_0_subtile_53__pin_clk_7_, bottom_width_0_height_0_subtile_53__pin_clk_8_, bottom_width_0_height_0_subtile_53__pin_clk_9_, bottom_width_0_height_0_subtile_53__pin_clk_10_, bottom_width_0_height_0_subtile_53__pin_clk_11_, bottom_width_0_height_0_subtile_53__pin_clk_12_, bottom_width_0_height_0_subtile_53__pin_clk_13_, bottom_width_0_height_0_subtile_53__pin_clk_14_, bottom_width_0_height_0_subtile_53__pin_clk_15_}),
		.ccff_head(logical_tile_io_corner_mode_io_corner__52_ccff_tail),
		.io_corner_a2f_o({top_width_0_height_0_subtile_53__pin_a2f_o_0_, top_width_0_height_0_subtile_53__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_53__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_corner_mode_io_corner__53_ccff_tail));

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__54 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[54]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[54]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[54]),
		.io_corner_f2a_i(top_width_0_height_0_subtile_54__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_54__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_54__pin_clk_0_, bottom_width_0_height_0_subtile_54__pin_clk_1_, bottom_width_0_height_0_subtile_54__pin_clk_2_, bottom_width_0_height_0_subtile_54__pin_clk_3_, bottom_width_0_height_0_subtile_54__pin_clk_4_, bottom_width_0_height_0_subtile_54__pin_clk_5_, bottom_width_0_height_0_subtile_54__pin_clk_6_, bottom_width_0_height_0_subtile_54__pin_clk_7_, bottom_width_0_height_0_subtile_54__pin_clk_8_, bottom_width_0_height_0_subtile_54__pin_clk_9_, bottom_width_0_height_0_subtile_54__pin_clk_10_, bottom_width_0_height_0_subtile_54__pin_clk_11_, bottom_width_0_height_0_subtile_54__pin_clk_12_, bottom_width_0_height_0_subtile_54__pin_clk_13_, bottom_width_0_height_0_subtile_54__pin_clk_14_, bottom_width_0_height_0_subtile_54__pin_clk_15_}),
		.ccff_head(logical_tile_io_corner_mode_io_corner__53_ccff_tail),
		.io_corner_a2f_o({top_width_0_height_0_subtile_54__pin_a2f_o_0_, top_width_0_height_0_subtile_54__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_54__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_corner_mode_io_corner__54_ccff_tail));

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__55 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[55]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[55]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[55]),
		.io_corner_f2a_i(top_width_0_height_0_subtile_55__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_55__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_55__pin_clk_0_, bottom_width_0_height_0_subtile_55__pin_clk_1_, bottom_width_0_height_0_subtile_55__pin_clk_2_, bottom_width_0_height_0_subtile_55__pin_clk_3_, bottom_width_0_height_0_subtile_55__pin_clk_4_, bottom_width_0_height_0_subtile_55__pin_clk_5_, bottom_width_0_height_0_subtile_55__pin_clk_6_, bottom_width_0_height_0_subtile_55__pin_clk_7_, bottom_width_0_height_0_subtile_55__pin_clk_8_, bottom_width_0_height_0_subtile_55__pin_clk_9_, bottom_width_0_height_0_subtile_55__pin_clk_10_, bottom_width_0_height_0_subtile_55__pin_clk_11_, bottom_width_0_height_0_subtile_55__pin_clk_12_, bottom_width_0_height_0_subtile_55__pin_clk_13_, bottom_width_0_height_0_subtile_55__pin_clk_14_, bottom_width_0_height_0_subtile_55__pin_clk_15_}),
		.ccff_head(logical_tile_io_corner_mode_io_corner__54_ccff_tail),
		.io_corner_a2f_o({top_width_0_height_0_subtile_55__pin_a2f_o_0_, top_width_0_height_0_subtile_55__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_55__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_corner_mode_io_corner__55_ccff_tail));

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__56 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[56]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[56]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[56]),
		.io_corner_f2a_i(top_width_0_height_0_subtile_56__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_56__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_56__pin_clk_0_, bottom_width_0_height_0_subtile_56__pin_clk_1_, bottom_width_0_height_0_subtile_56__pin_clk_2_, bottom_width_0_height_0_subtile_56__pin_clk_3_, bottom_width_0_height_0_subtile_56__pin_clk_4_, bottom_width_0_height_0_subtile_56__pin_clk_5_, bottom_width_0_height_0_subtile_56__pin_clk_6_, bottom_width_0_height_0_subtile_56__pin_clk_7_, bottom_width_0_height_0_subtile_56__pin_clk_8_, bottom_width_0_height_0_subtile_56__pin_clk_9_, bottom_width_0_height_0_subtile_56__pin_clk_10_, bottom_width_0_height_0_subtile_56__pin_clk_11_, bottom_width_0_height_0_subtile_56__pin_clk_12_, bottom_width_0_height_0_subtile_56__pin_clk_13_, bottom_width_0_height_0_subtile_56__pin_clk_14_, bottom_width_0_height_0_subtile_56__pin_clk_15_}),
		.ccff_head(logical_tile_io_corner_mode_io_corner__55_ccff_tail),
		.io_corner_a2f_o({top_width_0_height_0_subtile_56__pin_a2f_o_0_, top_width_0_height_0_subtile_56__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_56__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_corner_mode_io_corner__56_ccff_tail));

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__57 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[57]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[57]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[57]),
		.io_corner_f2a_i(top_width_0_height_0_subtile_57__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_57__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_57__pin_clk_0_, bottom_width_0_height_0_subtile_57__pin_clk_1_, bottom_width_0_height_0_subtile_57__pin_clk_2_, bottom_width_0_height_0_subtile_57__pin_clk_3_, bottom_width_0_height_0_subtile_57__pin_clk_4_, bottom_width_0_height_0_subtile_57__pin_clk_5_, bottom_width_0_height_0_subtile_57__pin_clk_6_, bottom_width_0_height_0_subtile_57__pin_clk_7_, bottom_width_0_height_0_subtile_57__pin_clk_8_, bottom_width_0_height_0_subtile_57__pin_clk_9_, bottom_width_0_height_0_subtile_57__pin_clk_10_, bottom_width_0_height_0_subtile_57__pin_clk_11_, bottom_width_0_height_0_subtile_57__pin_clk_12_, bottom_width_0_height_0_subtile_57__pin_clk_13_, bottom_width_0_height_0_subtile_57__pin_clk_14_, bottom_width_0_height_0_subtile_57__pin_clk_15_}),
		.ccff_head(logical_tile_io_corner_mode_io_corner__56_ccff_tail),
		.io_corner_a2f_o({top_width_0_height_0_subtile_57__pin_a2f_o_0_, top_width_0_height_0_subtile_57__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_57__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_corner_mode_io_corner__57_ccff_tail));

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__58 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[58]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[58]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[58]),
		.io_corner_f2a_i(top_width_0_height_0_subtile_58__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_58__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_58__pin_clk_0_, bottom_width_0_height_0_subtile_58__pin_clk_1_, bottom_width_0_height_0_subtile_58__pin_clk_2_, bottom_width_0_height_0_subtile_58__pin_clk_3_, bottom_width_0_height_0_subtile_58__pin_clk_4_, bottom_width_0_height_0_subtile_58__pin_clk_5_, bottom_width_0_height_0_subtile_58__pin_clk_6_, bottom_width_0_height_0_subtile_58__pin_clk_7_, bottom_width_0_height_0_subtile_58__pin_clk_8_, bottom_width_0_height_0_subtile_58__pin_clk_9_, bottom_width_0_height_0_subtile_58__pin_clk_10_, bottom_width_0_height_0_subtile_58__pin_clk_11_, bottom_width_0_height_0_subtile_58__pin_clk_12_, bottom_width_0_height_0_subtile_58__pin_clk_13_, bottom_width_0_height_0_subtile_58__pin_clk_14_, bottom_width_0_height_0_subtile_58__pin_clk_15_}),
		.ccff_head(logical_tile_io_corner_mode_io_corner__57_ccff_tail),
		.io_corner_a2f_o({top_width_0_height_0_subtile_58__pin_a2f_o_0_, top_width_0_height_0_subtile_58__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_58__pin_sc_out_0_),
		.ccff_tail(logical_tile_io_corner_mode_io_corner__58_ccff_tail));

	logical_tile_io_corner_mode_io_corner_ logical_tile_io_corner_mode_io_corner__59 (
		.global_reset(global_reset),
		.scan_mode(scan_mode),
		.scan_enable(scan_enable),
		.config_enable(config_enable),
		.prog_clock(prog_clock),
		.gfpga_pad_RS_PREIO_A2F(gfpga_pad_RS_PREIO_A2F[59]),
		.gfpga_pad_RS_PREIO_F2A(gfpga_pad_RS_PREIO_F2A[59]),
		.gfpga_pad_RS_PREIO_SOC_CLK(gfpga_pad_RS_PREIO_SOC_CLK[59]),
		.io_corner_f2a_i(top_width_0_height_0_subtile_59__pin_f2a_i_0_),
		.io_corner_sc_in(left_width_0_height_0_subtile_59__pin_sc_in_0_),
		.io_corner_clk({bottom_width_0_height_0_subtile_59__pin_clk_0_, bottom_width_0_height_0_subtile_59__pin_clk_1_, bottom_width_0_height_0_subtile_59__pin_clk_2_, bottom_width_0_height_0_subtile_59__pin_clk_3_, bottom_width_0_height_0_subtile_59__pin_clk_4_, bottom_width_0_height_0_subtile_59__pin_clk_5_, bottom_width_0_height_0_subtile_59__pin_clk_6_, bottom_width_0_height_0_subtile_59__pin_clk_7_, bottom_width_0_height_0_subtile_59__pin_clk_8_, bottom_width_0_height_0_subtile_59__pin_clk_9_, bottom_width_0_height_0_subtile_59__pin_clk_10_, bottom_width_0_height_0_subtile_59__pin_clk_11_, bottom_width_0_height_0_subtile_59__pin_clk_12_, bottom_width_0_height_0_subtile_59__pin_clk_13_, bottom_width_0_height_0_subtile_59__pin_clk_14_, bottom_width_0_height_0_subtile_59__pin_clk_15_}),
		.ccff_head(logical_tile_io_corner_mode_io_corner__58_ccff_tail),
		.io_corner_a2f_o({top_width_0_height_0_subtile_59__pin_a2f_o_0_, top_width_0_height_0_subtile_59__pin_a2f_o_1_}),
		.io_corner_sc_out(left_width_0_height_0_subtile_59__pin_sc_out_0_),
		.ccff_tail(ccff_tail));

endmodule
// ----- END Verilog module for grid_io_right_top -----

//----- Default net type -----
`default_nettype none



// ----- END Grid Verilog module: grid_io_right_top -----

