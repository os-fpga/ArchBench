//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for primitive pb_type: logic0
//	Author: Xifan TANG
//	Organization: University of Utah
//-------------------------------------------
//----- Time scale -----
`timescale 1ns / 1ps

//----- Default net type -----
`default_nettype wire

// ----- Verilog module for logical_tile_dsp_mode_default__opt_mode_default__logic0 -----
module logical_tile_dsp_mode_default__opt_mode_default__logic0(logic0_logic0);
//----- OUTPUT PORTS -----
output [0:0] logic0_logic0;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	logic0 logic0_0_ (
		.logic0(logic0_logic0));

endmodule
// ----- END Verilog module for logical_tile_dsp_mode_default__opt_mode_default__logic0 -----

//----- Default net type -----
`default_nettype none



